netcdf ostia_seaice_obs.cdl {
dimensions:
	nlocs = 11 ;
	nvars = 1 ;
	ndatetime = 20 ;
	nstring = 50 ;
variables:
	float ndatetime(ndatetime) ;
		ndatetime:suggested_chunk_dim = 100LL ;
	float nlocs(nlocs) ;
		nlocs:suggested_chunk_dim = 100LL ;
	float nstring(nstring) ;
		nstring:suggested_chunk_dim = 100LL ;
	float nvars(nvars) ;
		nvars:suggested_chunk_dim = 100LL ;

// global attributes:
		string :_ioda_layout = "ObsGroup" ;
		:_ioda_layout_version = 0 ;
		:nvars = 1 ;
		:date_time = 2021070100 ;
		:odb_version = 2LL ;
		:history = "Mon Aug 23 11:00:30 2021: ncks --fix_rec_dmn nlocs tmp2.nc obs_seaice_20210701T0000Z_v_reduced.nc4\nMon Aug 23 11:00:20 2021: ncrcat -d nlocs,1,,1000000 tmp.nc tmp2.nc\nSat Aug 21 17:00:19 2021: ncks --mk_rec_dmn nlocs obs_seaice_20210701T0000Z.nc4 tmp.nc" ;
		:NCO = "netCDF Operators version 4.7.5 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
		:nco_openmp_thread_number = 1 ;
		:nlocs = 11 ;
data:

 ndatetime = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 nlocs = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 nstring = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0 ;

 nvars = 0 ;

group: MetaData {
  variables:
  	string datetime(nlocs) ;
  	float latitude(nlocs) ;
  	float longitude(nlocs) ;
  	int ops_obsgroup(nlocs) ;
  	int ops_subtype(nlocs) ;
  	int record_number(nlocs) ;
  	int sequence_number(nlocs) ;
  	float time(nlocs) ;
  data:

   datetime = "2021-06-29T12:00:00Z", "2021-06-29T12:00:00Z", 
      "2021-06-29T12:00:00Z", "2021-06-29T12:00:00Z", "2021-06-30T00:00:00Z", 
      "2021-06-30T00:00:00Z", "2021-06-30T00:00:00Z", "2021-06-30T00:00:00Z", 
      "2021-06-30T00:00:00Z", "2021-06-30T00:00:00Z", "2021-06-30T00:00:00Z" ;

   latitude = 82.02939, 62.43589, -65.28536, -51.87979, 41.8942, 22.6519, 
      3.3263, -15.916, -35.2416, -54.4839, -73.7262 ;

   longitude = 168.338, 31.21495, -24.91501, -154.482, 38.443, -148.293, 
      25.115, -161.621, 11.787, -174.949, -1.685 ;

   ops_obsgroup = 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30 ;

   ops_subtype = 60700, 60700, 60700, 60700, 60600, 60600, 60600, 60600, 
      60600, 60600, 60600 ;

   record_number = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

   sequence_number = 1, 500001, 1000001, 1500001, 2493102, 3493102, 4493102, 
      5493102, 6493102, 7493102, 8493102 ;

   time = -12, -12, -12, -12, -24, -24, -24, -24, -24, -24, -24 ;
  } // group MetaData

group: ObsError {
  variables:
  	float ice_area_fraction(nlocs) ;
  data:

   ice_area_fraction = 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1 ;
  } // group ObsError

group: ObsValue {
  variables:
  	float ice_area_fraction(nlocs) ;
  data:

   ice_area_fraction = 0, _, 0.9963, 0, 0, 0, 0, 0, 0, 0, 0 ;
  } // group ObsValue

group: PreQC {
  variables:
  	float ice_area_fraction(nlocs) ;
  data:

   ice_area_fraction = 1e+09, 1e+09, 1e+09, 1e+09, 1e+09, 1e+09, 1e+09, 
      1e+09, 1e+09, 1e+09, 1e+09 ;
  } // group PreQC

group: VarMetaData {
  variables:
  	string variable_names(nvars) ;
  data:

   variable_names = "ice_area_fraction" ;
  } // group VarMetaData
}
