netcdf simple_fdbk {
dimensions:
	x = 3 ;
	y = 2 ;
        t = 1 ; 
variables:
        double nav_lat(y, x) ;
	double nav_lon(y, x) ;
        double iiceconc(t, y, x) ;
        int t(t);
            t:units = "seconds since 1970-01-01 00:00:00" ;

data:

 t = 0;

 nav_lat =
  0, 0, 0,
  1, 1, 1;
 
 nav_lon =
  10, 11, 12,
  10, 11, 12;

 iiceconc =
  120, 130, 140,
  150, 160, 170;
}
