netcdf simple_fdbk {
dimensions:
	x = 3 ;
	y = 2 ;
        t = 3 ;
variables:
        double nav_lat(y, x) ;
	double nav_lon(y, x) ;
        double iiceconc(t, y, x) ;
            iiceconc:_FillValue = -32768 ;
        int t(t);
            t:units = "seconds since 1970-01-01 00:00:00" ;

data:

 t = 0, 86400, 172800;

 nav_lat =
  0, 0, 0,
  1, 1, 1;

 nav_lon =
  10, 11, 12,
  10, 11, 12;

 iiceconc =
  120, 130, 140,
  150, 160, 170,
  121, 131, 141,
  151, 161, 171,
  122, 132, 142,
  152, 162, 172 ;

}
