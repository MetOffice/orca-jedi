netcdf orca2_t_bkg {
dimensions:
	x = 182 ;
	y = 149 ;
	z = 2 ;
	t = 1 ;
variables:
	double nav_lat(y, x) ;
	double nav_lon(y, x) ;
        int t(t) ;
            t:units = "seconds since 1981-01-01 00:00:00" ;
	double sic_tot_var(t, y, x) ;
data:

 t = 0;

 nav_lat =
  -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, 
    -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, 
    -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, 
    -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, 
    -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, 
    -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, 
    -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, 
    -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, 
    -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, 
    -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, 
    -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, 
    -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, 
    -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, 
    -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, 
    -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, 
    -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, 
    -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, 
    -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, 
    -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, 
    -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, 
    -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, 
    -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, 
    -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, 
    -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, 
    -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, 
    -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, 
    -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, 
    -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, 
    -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, 
    -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, -78.19058, 
    -78.19058, -78.19058,
  -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, 
    -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, 
    -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, 
    -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, 
    -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, 
    -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, 
    -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, 
    -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, 
    -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, 
    -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, 
    -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, 
    -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, 
    -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, 
    -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, 
    -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, 
    -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, 
    -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, 
    -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, 
    -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, 
    -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, 
    -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, 
    -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, 
    -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, 
    -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, 
    -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, 
    -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742, -77.7742,
  -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, 
    -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, 
    -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, 
    -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, 
    -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, 
    -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, 
    -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, 
    -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, 
    -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, 
    -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, 
    -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, 
    -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, 
    -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, 
    -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, 
    -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, 
    -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, 
    -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, 
    -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, 
    -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, 
    -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, 
    -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, 
    -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, 
    -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, 
    -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, 
    -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, 
    -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, 
    -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, 
    -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, 
    -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, 
    -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, -77.34337, 
    -77.34337, -77.34337,
  -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, 
    -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, 
    -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, 
    -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, 
    -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, 
    -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, 
    -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, 
    -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, 
    -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, 
    -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, 
    -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, 
    -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, 
    -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, 
    -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, 
    -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, 
    -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, 
    -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, 
    -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, 
    -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, 
    -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, 
    -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, 
    -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, 
    -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, 
    -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, 
    -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, 
    -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, 
    -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, 
    -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, 
    -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, 
    -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, -76.89761, 
    -76.89761, -76.89761,
  -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, 
    -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, 
    -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, 
    -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, 
    -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, 
    -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, 
    -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, 
    -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, 
    -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, 
    -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, 
    -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, 
    -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, 
    -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, 
    -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, 
    -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, 
    -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, 
    -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, 
    -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, 
    -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, 
    -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, 
    -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, 
    -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, 
    -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, 
    -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, 
    -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, 
    -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, 
    -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, 
    -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, 
    -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, 
    -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, -76.43644, 
    -76.43644, -76.43644,
  -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, 
    -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, 
    -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, 
    -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, 
    -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, 
    -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, 
    -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, 
    -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, 
    -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, 
    -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, 
    -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, 
    -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, 
    -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, 
    -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, 
    -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, 
    -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, 
    -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, 
    -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, 
    -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, 
    -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, 
    -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, 
    -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, 
    -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, 
    -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, 
    -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, 
    -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, 
    -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, 
    -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, 
    -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, 
    -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, -75.95934, 
    -75.95934, -75.95934,
  -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, 
    -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, 
    -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, 
    -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, 
    -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, 
    -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, 
    -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, 
    -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, 
    -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, 
    -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, 
    -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, 
    -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, 
    -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, 
    -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, 
    -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, 
    -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, 
    -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, 
    -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, 
    -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, 
    -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, 
    -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, 
    -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, 
    -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, 
    -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, 
    -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, 
    -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, 
    -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, 
    -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, 
    -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, 
    -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, -75.46582, 
    -75.46582, -75.46582,
  -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, 
    -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, 
    -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, 
    -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, 
    -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, 
    -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, 
    -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, 
    -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, 
    -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, 
    -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, 
    -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, 
    -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, 
    -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, 
    -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, 
    -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, 
    -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, 
    -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, 
    -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, 
    -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, 
    -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, 
    -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, 
    -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, 
    -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, 
    -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, 
    -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, 
    -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, 
    -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, 
    -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, 
    -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, 
    -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, -74.95534, 
    -74.95534, -74.95534,
  -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, 
    -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, 
    -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, 
    -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, 
    -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, 
    -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, 
    -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, 
    -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, 
    -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, 
    -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, 
    -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, 
    -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, 
    -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, 
    -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, 
    -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, 
    -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, 
    -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, 
    -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, 
    -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, 
    -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, 
    -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, 
    -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, 
    -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, 
    -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, 
    -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, 
    -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, 
    -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, 
    -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, 
    -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, 
    -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, -74.42735, 
    -74.42735, -74.42735,
  -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, 
    -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, 
    -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, 
    -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, 
    -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, 
    -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, 
    -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, 
    -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, 
    -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, 
    -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, 
    -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, 
    -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, 
    -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, 
    -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, 
    -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, 
    -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, 
    -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, 
    -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, 
    -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, 
    -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, 
    -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, 
    -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, 
    -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, 
    -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, 
    -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, 
    -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, 
    -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, 
    -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, 
    -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, 
    -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, -73.88131, 
    -73.88131, -73.88131,
  -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, 
    -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, 
    -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, 
    -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, 
    -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, 
    -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, 
    -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, 
    -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, 
    -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, 
    -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, 
    -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, 
    -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, 
    -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, 
    -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, 
    -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, 
    -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, 
    -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, 
    -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, 
    -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, 
    -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, 
    -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, 
    -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, 
    -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, 
    -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, 
    -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, 
    -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, 
    -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, 
    -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, 
    -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, 
    -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, -73.31665, 
    -73.31665, -73.31665,
  -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, 
    -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, 
    -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, 
    -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, 
    -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, 
    -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, 
    -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, 
    -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, 
    -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, 
    -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, 
    -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, 
    -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, 
    -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, 
    -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, 
    -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, 
    -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, 
    -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, 
    -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, 
    -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, 
    -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, 
    -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, 
    -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, 
    -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, 
    -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, 
    -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, 
    -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, 
    -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, 
    -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, 
    -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, 
    -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, -72.73279, 
    -72.73279, -72.73279,
  -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, 
    -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, 
    -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, 
    -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, 
    -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, 
    -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, 
    -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, 
    -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, 
    -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, 
    -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, 
    -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, 
    -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, 
    -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, 
    -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, 
    -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, 
    -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, 
    -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, 
    -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, 
    -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, 
    -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, 
    -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, 
    -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, 
    -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, 
    -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, 
    -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, 
    -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, 
    -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, 
    -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, 
    -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, 
    -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, -72.12914, 
    -72.12914, -72.12914,
  -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, 
    -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, 
    -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, 
    -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, 
    -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, 
    -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, 
    -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, 
    -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, 
    -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, 
    -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, 
    -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, 
    -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, 
    -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, 
    -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, 
    -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, 
    -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, 
    -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, 
    -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, 
    -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, 
    -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, 
    -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, 
    -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, 
    -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, 
    -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, 
    -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, 
    -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051, -71.5051,
  -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, 
    -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, 
    -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, 
    -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, 
    -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, 
    -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, 
    -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, 
    -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, 
    -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, 
    -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, 
    -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, 
    -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, 
    -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, 
    -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, 
    -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, 
    -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, 
    -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, 
    -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, 
    -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, 
    -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, 
    -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, 
    -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, 
    -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, 
    -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, 
    -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, 
    -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, 
    -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, 
    -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, 
    -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, 
    -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, -70.86005, 
    -70.86005, -70.86005,
  -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, 
    -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, 
    -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, 
    -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, 
    -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, 
    -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, 
    -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, 
    -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, 
    -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, 
    -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, 
    -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, 
    -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, 
    -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, 
    -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, 
    -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, 
    -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, 
    -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, 
    -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, 
    -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, 
    -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, 
    -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, 
    -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, 
    -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, 
    -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, 
    -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, 
    -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, 
    -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, 
    -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, 
    -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, 
    -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, -70.19337, 
    -70.19337, -70.19337,
  -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, 
    -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, 
    -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, 
    -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, 
    -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, 
    -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, 
    -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, 
    -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, 
    -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, 
    -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, 
    -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, 
    -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, 
    -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, 
    -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, 
    -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, 
    -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, 
    -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, 
    -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, 
    -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, 
    -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, 
    -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, 
    -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, 
    -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, 
    -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, 
    -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, 
    -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, 
    -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, 
    -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, 
    -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, 
    -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, -69.50445, 
    -69.50445, -69.50445,
  -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, 
    -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, 
    -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, 
    -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, 
    -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, 
    -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, 
    -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, 
    -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, 
    -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, 
    -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, 
    -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, 
    -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, 
    -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, 
    -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, 
    -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, 
    -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, 
    -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, 
    -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, 
    -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, 
    -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, 
    -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, 
    -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, 
    -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, 
    -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, 
    -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, 
    -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, 
    -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, 
    -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, 
    -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, 
    -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, -68.79263, 
    -68.79263, -68.79263,
  -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, 
    -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, 
    -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, 
    -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, 
    -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, 
    -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, 
    -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, 
    -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, 
    -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, 
    -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, 
    -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, 
    -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, 
    -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, 
    -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, 
    -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, 
    -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, 
    -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, 
    -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, 
    -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, 
    -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, 
    -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, 
    -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, 
    -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, 
    -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, 
    -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, 
    -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, 
    -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, 
    -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, 
    -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, 
    -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, -68.05725, 
    -68.05725, -68.05725,
  -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, 
    -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, 
    -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, 
    -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, 
    -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, 
    -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, 
    -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, 
    -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, 
    -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, 
    -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, 
    -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, 
    -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, 
    -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, 
    -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, 
    -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, 
    -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, 
    -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, 
    -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, 
    -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, 
    -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, 
    -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, 
    -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, 
    -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, 
    -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, 
    -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, 
    -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, 
    -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, 
    -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, 
    -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, 
    -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, -67.29768, 
    -67.29768, -67.29768,
  -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, 
    -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, 
    -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, 
    -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, 
    -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, 
    -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, 
    -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, 
    -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, 
    -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, 
    -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, 
    -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, 
    -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, 
    -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, 
    -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, 
    -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, 
    -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, 
    -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, 
    -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, 
    -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, 
    -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, 
    -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, 
    -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, 
    -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, 
    -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, 
    -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, 
    -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, 
    -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, 
    -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, 
    -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, 
    -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, -66.51326, 
    -66.51326, -66.51326,
  -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, 
    -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, 
    -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, 
    -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, 
    -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, 
    -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, 
    -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, 
    -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, 
    -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, 
    -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, 
    -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, 
    -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, 
    -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, 
    -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, 
    -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, 
    -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, 
    -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, 
    -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, 
    -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, 
    -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, 
    -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, 
    -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, 
    -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, 
    -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, 
    -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, 
    -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, 
    -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, 
    -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, 
    -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, 
    -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, -65.70332, 
    -65.70332, -65.70332,
  -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, 
    -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, 
    -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, 
    -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, 
    -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, 
    -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, 
    -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, 
    -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, 
    -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, 
    -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, 
    -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, 
    -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, 
    -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, 
    -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, 
    -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, 
    -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, 
    -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, 
    -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, 
    -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, 
    -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, 
    -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, 
    -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, 
    -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, 
    -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, 
    -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, 
    -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672, -64.8672,
  -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, 
    -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, 
    -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, 
    -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, 
    -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, 
    -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, 
    -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, 
    -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, 
    -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, 
    -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, 
    -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, 
    -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, 
    -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, 
    -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, 
    -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, 
    -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, 
    -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, 
    -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, 
    -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, 
    -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, 
    -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, 
    -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, 
    -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, 
    -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, 
    -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, 
    -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, 
    -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, 
    -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, 
    -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, 
    -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, -64.00423, 
    -64.00423, -64.00423,
  -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, 
    -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, 
    -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, 
    -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, 
    -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, 
    -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, 
    -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, 
    -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, 
    -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, 
    -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, 
    -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, 
    -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, 
    -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, 
    -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, 
    -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, 
    -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, 
    -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, 
    -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, 
    -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, 
    -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, 
    -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, 
    -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, 
    -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, 
    -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, 
    -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, 
    -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, 
    -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, 
    -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, 
    -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, 
    -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, -63.11375, 
    -63.11375, -63.11375,
  -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, 
    -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, 
    -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, 
    -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, 
    -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, 
    -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, 
    -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, 
    -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, 
    -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, 
    -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, 
    -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, 
    -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, 
    -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, 
    -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, 
    -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, 
    -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, 
    -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, 
    -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, 
    -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, 
    -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, 
    -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, 
    -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, 
    -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, 
    -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, 
    -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, 
    -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, 
    -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, 
    -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, 
    -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, 
    -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, -62.19513, 
    -62.19513, -62.19513,
  -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, 
    -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, 
    -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, 
    -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, 
    -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, 
    -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, 
    -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, 
    -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, 
    -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, 
    -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, 
    -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, 
    -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, 
    -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, 
    -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, 
    -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, 
    -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, 
    -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, 
    -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, 
    -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, 
    -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, 
    -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, 
    -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, 
    -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, 
    -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, 
    -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, 
    -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, 
    -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, 
    -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, 
    -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, 
    -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, -61.24769, 
    -61.24769, -61.24769,
  -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, 
    -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, 
    -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, 
    -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, 
    -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, 
    -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, 
    -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, 
    -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, 
    -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, 
    -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, 
    -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, 
    -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, 
    -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, 
    -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, 
    -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, 
    -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, 
    -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, 
    -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, 
    -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, 
    -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, 
    -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, 
    -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, 
    -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, 
    -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, 
    -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, 
    -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, 
    -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, 
    -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, 
    -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, 
    -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, -60.27082, 
    -60.27082, -60.27082,
  -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, 
    -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, 
    -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, 
    -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, 
    -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, 
    -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, 
    -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, 
    -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, 
    -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, 
    -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, 
    -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, 
    -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, 
    -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, 
    -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, 
    -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, 
    -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, 
    -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, 
    -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, 
    -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, 
    -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, 
    -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, 
    -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, 
    -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, 
    -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, 
    -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, 
    -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, 
    -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, 
    -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, 
    -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, 
    -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, -59.26389, 
    -59.26389, -59.26389,
  -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, 
    -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, 
    -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, 
    -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, 
    -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, 
    -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, 
    -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, 
    -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, 
    -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, 
    -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, 
    -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, 
    -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, 
    -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, 
    -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, 
    -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, 
    -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, 
    -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, 
    -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, 
    -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, 
    -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, 
    -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, 
    -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, 
    -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, 
    -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, 
    -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, 
    -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, 
    -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, 
    -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, 
    -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, 
    -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, -58.22628, 
    -58.22628, -58.22628,
  -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, 
    -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, 
    -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, 
    -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, 
    -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, 
    -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, 
    -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, 
    -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, 
    -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, 
    -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, 
    -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, 
    -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, 
    -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, 
    -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, 
    -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, 
    -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, 
    -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, 
    -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, 
    -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, 
    -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, 
    -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, 
    -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, 
    -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, 
    -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, 
    -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, 
    -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, 
    -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, 
    -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, 
    -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, 
    -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, -57.15743, 
    -57.15743, -57.15743,
  -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, 
    -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, 
    -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, 
    -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, 
    -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, 
    -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, 
    -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, 
    -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, 
    -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, 
    -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, 
    -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, 
    -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, 
    -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, 
    -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, 
    -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, 
    -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, 
    -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, 
    -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, 
    -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, 
    -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, 
    -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, 
    -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, 
    -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, 
    -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, 
    -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, 
    -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, 
    -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, 
    -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, 
    -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, 
    -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, -56.05677, 
    -56.05677, -56.05677,
  -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, 
    -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, 
    -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, 
    -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, 
    -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, 
    -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, 
    -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, 
    -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, 
    -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, 
    -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, 
    -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, 
    -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, 
    -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, 
    -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, 
    -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, 
    -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, 
    -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, 
    -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, 
    -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, 
    -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, 
    -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, 
    -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, 
    -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, 
    -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, 
    -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, 
    -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, 
    -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, 
    -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, 
    -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, 
    -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, -54.92377, 
    -54.92377, -54.92377,
  -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, 
    -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, 
    -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, 
    -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, 
    -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, 
    -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, 
    -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, 
    -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, 
    -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, 
    -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, 
    -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, 
    -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, 
    -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, 
    -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, 
    -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, 
    -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, 
    -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, 
    -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, 
    -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, 
    -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, 
    -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, 
    -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, 
    -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, 
    -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, 
    -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, 
    -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, 
    -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, 
    -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, 
    -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, 
    -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, -53.75795, 
    -53.75795, -53.75795,
  -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, 
    -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, 
    -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, 
    -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, 
    -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, 
    -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, 
    -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, 
    -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, 
    -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, 
    -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, 
    -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, 
    -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, 
    -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, 
    -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, 
    -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, 
    -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, 
    -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, 
    -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, 
    -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, 
    -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, 
    -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, 
    -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, 
    -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, 
    -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, 
    -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, 
    -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, 
    -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, 
    -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, 
    -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, 
    -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, -52.55884, 
    -52.55884, -52.55884,
  -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, 
    -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, 
    -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, 
    -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, 
    -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, 
    -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, 
    -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, 
    -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, 
    -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, 
    -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, 
    -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, 
    -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, 
    -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, 
    -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, 
    -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, 
    -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, 
    -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, 
    -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, 
    -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, 
    -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, 
    -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, 
    -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, 
    -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, 
    -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, 
    -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, 
    -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, 
    -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, 
    -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, 
    -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, 
    -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, -51.32603, 
    -51.32603, -51.32603,
  -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, 
    -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, 
    -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, 
    -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, 
    -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, 
    -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, 
    -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, 
    -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, 
    -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, 
    -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, 
    -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, 
    -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, 
    -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, 
    -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, 
    -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, 
    -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, 
    -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, 
    -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, 
    -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, 
    -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, 
    -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, 
    -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, 
    -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, 
    -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, 
    -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, 
    -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, 
    -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, 
    -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, 
    -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, 
    -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, -50.05918, 
    -50.05918, -50.05918,
  -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, 
    -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, 
    -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, 
    -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, 
    -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, 
    -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, 
    -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, 
    -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, 
    -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, 
    -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, 
    -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, 
    -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, 
    -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, 
    -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, 
    -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, 
    -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, 
    -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, 
    -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, 
    -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, 
    -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, 
    -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, 
    -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, 
    -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, 
    -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, 
    -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, 
    -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, 
    -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, 
    -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, 
    -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, 
    -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, -48.75796, 
    -48.75796, -48.75796,
  -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, 
    -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, 
    -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, 
    -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, 
    -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, 
    -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, 
    -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, 
    -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, 
    -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, 
    -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, 
    -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, 
    -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, 
    -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, 
    -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, 
    -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, 
    -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, 
    -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, 
    -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, 
    -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, 
    -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, 
    -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, 
    -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, 
    -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, 
    -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, 
    -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, 
    -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, 
    -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, 
    -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, 
    -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, 
    -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, -47.42214, 
    -47.42214, -47.42214,
  -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, 
    -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, 
    -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, 
    -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, 
    -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, 
    -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, 
    -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, 
    -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, 
    -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, 
    -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, 
    -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, 
    -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, 
    -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, 
    -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, 
    -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, 
    -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, 
    -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, 
    -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, 
    -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, 
    -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, 
    -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, 
    -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, 
    -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, 
    -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, 
    -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, 
    -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, 
    -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, 
    -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, 
    -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, 
    -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, -46.05155, 
    -46.05155, -46.05155,
  -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, 
    -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, 
    -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, 
    -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, 
    -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, 
    -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, 
    -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, 
    -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, 
    -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, 
    -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, 
    -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, 
    -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, 
    -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, 
    -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, 
    -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, 
    -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, 
    -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, 
    -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, 
    -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, 
    -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, 
    -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, 
    -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, 
    -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, 
    -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, 
    -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, 
    -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, 
    -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, 
    -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, 
    -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, 
    -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, -44.64608, 
    -44.64608, -44.64608,
  -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, 
    -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, 
    -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, 
    -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, 
    -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, 
    -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, 
    -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, 
    -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, 
    -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, 
    -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, 
    -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, 
    -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, 
    -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, 
    -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, 
    -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, 
    -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, 
    -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, 
    -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, 
    -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, 
    -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, 
    -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, 
    -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, 
    -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, 
    -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, 
    -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, 
    -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, 
    -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, 
    -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, 
    -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, 
    -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, -43.20571, 
    -43.20571, -43.20571,
  -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, 
    -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, 
    -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, 
    -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, 
    -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, 
    -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, 
    -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, 
    -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, 
    -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, 
    -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, 
    -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, 
    -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, 
    -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, 
    -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, 
    -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, 
    -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, 
    -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, 
    -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, 
    -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, 
    -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, 
    -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, 
    -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, 
    -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, 
    -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, 
    -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, 
    -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, 
    -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, 
    -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, 
    -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, 
    -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, -41.73051, 
    -41.73051, -41.73051,
  -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, 
    -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, 
    -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, 
    -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, 
    -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, 
    -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, 
    -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, 
    -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, 
    -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, 
    -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, 
    -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, 
    -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, 
    -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, 
    -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, 
    -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, 
    -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, 
    -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, 
    -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, 
    -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, 
    -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, 
    -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, 
    -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, 
    -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, 
    -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, 
    -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, 
    -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, 
    -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, 
    -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, 
    -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, 
    -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, -40.22064, 
    -40.22064, -40.22064,
  -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, 
    -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, 
    -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, 
    -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, 
    -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, 
    -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, 
    -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, 
    -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, 
    -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, 
    -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, 
    -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, 
    -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, 
    -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, 
    -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, 
    -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, 
    -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, 
    -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, 
    -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, 
    -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, 
    -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, 
    -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, 
    -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, 
    -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, 
    -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, 
    -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, 
    -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, 
    -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, 
    -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, 
    -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, 
    -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, -38.67636, 
    -38.67636, -38.67636,
  -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, 
    -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, 
    -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, 
    -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, 
    -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, 
    -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, 
    -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, 
    -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, 
    -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, 
    -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, 
    -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, 
    -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, 
    -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, 
    -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, 
    -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, 
    -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, 
    -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, 
    -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, 
    -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, 
    -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, 
    -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, 
    -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, 
    -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, 
    -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, 
    -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, 
    -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, 
    -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, 
    -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, 
    -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, 
    -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, -37.09803, 
    -37.09803, -37.09803,
  -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, 
    -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, 
    -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, 
    -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, 
    -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, 
    -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, 
    -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, 
    -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, 
    -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, 
    -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, 
    -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, 
    -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, 
    -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, 
    -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, 
    -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, 
    -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, 
    -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, 
    -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, 
    -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, 
    -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, 
    -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, 
    -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, 
    -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, 
    -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, 
    -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, 
    -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, 
    -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, 
    -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, 
    -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, 
    -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, -35.48612, 
    -35.48612, -35.48612,
  -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, 
    -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, 
    -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, 
    -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, 
    -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, 
    -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, 
    -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, 
    -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, 
    -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, 
    -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, 
    -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, 
    -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, 
    -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, 
    -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, 
    -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, 
    -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, 
    -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, 
    -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, 
    -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, 
    -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, 
    -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, 
    -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, 
    -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, 
    -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, 
    -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, 
    -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, 
    -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, 
    -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, 
    -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, 
    -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, -33.84122, 
    -33.84122, -33.84122,
  -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, 
    -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, 
    -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, 
    -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, 
    -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, 
    -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, 
    -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, 
    -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, 
    -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, 
    -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, 
    -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, 
    -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, 
    -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, 
    -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, 
    -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, 
    -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, 
    -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, 
    -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, 
    -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, 
    -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, 
    -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, 
    -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, 
    -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, 
    -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, 
    -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, 
    -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, 
    -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, 
    -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, 
    -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, 
    -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, -32.16404, 
    -32.16404, -32.16404,
  -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, 
    -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, 
    -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, 
    -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, 
    -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, 
    -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, 
    -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, 
    -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, 
    -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, 
    -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, 
    -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, 
    -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, 
    -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, 
    -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, 
    -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, 
    -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, 
    -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, 
    -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, 
    -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, 
    -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, 
    -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, 
    -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, 
    -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, 
    -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, 
    -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, 
    -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, 
    -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, 
    -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, 
    -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, 
    -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, -30.45541, 
    -30.45541, -30.45541,
  -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, 
    -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, 
    -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, 
    -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, 
    -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, 
    -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, 
    -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, 
    -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, 
    -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, 
    -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, 
    -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, 
    -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, 
    -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, 
    -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, 
    -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, 
    -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, 
    -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, 
    -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, 
    -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, 
    -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, 
    -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, 
    -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, 
    -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, 
    -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, 
    -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, 
    -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, 
    -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, 
    -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, 
    -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, 
    -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, -28.71628, 
    -28.71628, -28.71628,
  -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, 
    -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, 
    -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, 
    -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, 
    -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, 
    -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, 
    -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, 
    -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, 
    -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, 
    -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, 
    -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, 
    -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, 
    -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, 
    -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, 
    -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, 
    -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, 
    -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, 
    -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, 
    -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, 
    -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, 
    -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, 
    -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, 
    -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, 
    -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, 
    -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, 
    -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, 
    -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, 
    -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, 
    -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, 
    -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, -26.94775, 
    -26.94775, -26.94775,
  -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, 
    -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, 
    -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, 
    -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, 
    -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, 
    -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, 
    -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, 
    -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, 
    -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, 
    -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, 
    -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, 
    -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, 
    -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, 
    -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, 
    -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, 
    -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, 
    -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, 
    -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, 
    -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, 
    -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, 
    -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, 
    -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, 
    -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, 
    -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, 
    -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, 
    -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, 
    -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, 
    -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, 
    -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, 
    -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, -25.15103, 
    -25.15103, -25.15103,
  -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, 
    -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, 
    -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, 
    -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, 
    -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, 
    -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, 
    -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, 
    -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, 
    -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, 
    -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, 
    -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, 
    -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, 
    -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, 
    -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, 
    -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, 
    -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, 
    -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, 
    -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, 
    -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, 
    -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, 
    -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, 
    -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, 
    -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, 
    -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, 
    -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, 
    -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, 
    -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, 
    -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, 
    -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, 
    -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, -23.32746, 
    -23.32746, -23.32746,
  -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, 
    -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, 
    -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, 
    -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, 
    -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, 
    -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, 
    -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, 
    -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, 
    -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, 
    -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, 
    -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, 
    -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, 
    -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, 
    -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, 
    -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, 
    -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, 
    -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, 
    -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, 
    -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, 
    -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, 
    -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, 
    -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, 
    -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, 
    -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, 
    -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, 
    -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, 
    -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, 
    -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, 
    -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, 
    -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, -21.47852, 
    -21.47852, -21.47852,
  -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, 
    -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, 
    -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, 
    -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, 
    -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, 
    -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, 
    -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, 
    -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, 
    -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, 
    -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, 
    -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, 
    -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, 
    -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, 
    -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, 
    -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, 
    -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, 
    -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, 
    -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, 
    -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, 
    -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, 
    -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, 
    -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, 
    -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, 
    -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, 
    -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, 
    -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, 
    -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, 
    -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, 
    -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, 
    -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, -19.60579, 
    -19.60579, -19.60579,
  -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, 
    -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, 
    -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, 
    -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, 
    -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, 
    -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, 
    -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, 
    -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, 
    -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, 
    -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, 
    -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, 
    -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, 
    -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, 
    -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, 
    -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, 
    -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, 
    -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, 
    -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, 
    -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, 
    -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, 
    -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, 
    -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, 
    -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, 
    -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, 
    -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, 
    -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, 
    -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, 
    -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, 
    -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, 
    -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, -17.71952, 
    -17.71952, -17.71952,
  -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, 
    -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, 
    -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, 
    -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, 
    -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, 
    -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, 
    -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, 
    -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, 
    -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, 
    -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, 
    -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, 
    -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, 
    -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, 
    -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, 
    -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, 
    -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, 
    -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, 
    -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, 
    -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, 
    -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, 
    -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, 
    -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, 
    -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, 
    -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, 
    -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, 
    -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, 
    -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, 
    -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, 
    -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, 
    -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, -15.86032, 
    -15.86032, -15.86032,
  -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, 
    -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, 
    -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, 
    -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, 
    -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, 
    -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, 
    -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, 
    -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, 
    -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, 
    -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, 
    -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, 
    -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, 
    -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, 
    -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, 
    -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, 
    -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, 
    -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, 
    -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, 
    -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, 
    -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, 
    -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, 
    -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, 
    -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, 
    -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, 
    -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, 
    -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676, -14.0676,
  -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, 
    -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, 
    -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, 
    -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, 
    -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, 
    -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, 
    -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, 
    -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, 
    -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, 
    -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, 
    -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, 
    -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, 
    -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, 
    -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, 
    -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, 
    -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, 
    -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, 
    -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, 
    -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, 
    -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, 
    -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, 
    -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, 
    -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, 
    -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, 
    -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, 
    -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, 
    -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, 
    -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, 
    -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, 
    -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, -12.37097, 
    -12.37097, -12.37097,
  -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, 
    -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, 
    -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, 
    -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, 
    -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, 
    -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, 
    -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, 
    -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, 
    -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, 
    -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, 
    -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, 
    -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, 
    -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, 
    -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, 
    -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, 
    -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, 
    -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, 
    -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, 
    -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, 
    -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, 
    -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, 
    -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, 
    -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, 
    -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, 
    -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, 
    -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912, -10.7912,
  -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, 
    -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, 
    -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, 
    -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, 
    -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, 
    -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, 
    -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, 
    -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, 
    -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, 
    -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, 
    -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, 
    -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, 
    -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, 
    -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, 
    -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, 
    -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, 
    -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, 
    -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, 
    -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, 
    -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, 
    -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, 
    -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, 
    -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, 
    -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, 
    -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, 
    -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, 
    -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, 
    -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, 
    -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, 
    -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, -9.341137, 
    -9.341137, -9.341137,
  -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, 
    -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, 
    -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, 
    -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, 
    -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, 
    -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, 
    -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, 
    -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, 
    -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, 
    -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, 
    -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, 
    -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, 
    -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, 
    -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, 
    -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, 
    -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, 
    -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, 
    -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, 
    -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, 
    -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, 
    -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, 
    -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, 
    -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, 
    -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, 
    -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, 
    -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, 
    -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, 
    -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, 
    -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, 
    -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, -8.026655, 
    -8.026655, -8.026655,
  -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, 
    -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, 
    -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, 
    -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, 
    -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, 
    -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, 
    -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, 
    -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, 
    -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, 
    -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, 
    -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, 
    -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, 
    -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, 
    -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, 
    -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, 
    -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, 
    -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, 
    -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, 
    -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, 
    -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, 
    -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, 
    -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, 
    -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, 
    -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, 
    -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, 
    -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, 
    -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, 
    -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, 
    -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, 
    -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, -6.847561, 
    -6.847561, -6.847561,
  -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, 
    -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, 
    -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, 
    -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, 
    -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, 
    -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, 
    -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, 
    -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, 
    -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, 
    -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, 
    -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, 
    -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, 
    -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, 
    -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, 
    -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, 
    -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, 
    -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, 
    -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, 
    -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, 
    -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, 
    -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, 
    -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, 
    -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, 
    -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, 
    -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, 
    -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, 
    -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, 
    -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, 
    -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, 
    -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, -5.798548, 
    -5.798548, -5.798548,
  -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, 
    -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, 
    -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, 
    -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, 
    -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, 
    -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, 
    -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, 
    -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, 
    -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, 
    -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, 
    -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, 
    -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, 
    -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, 
    -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, 
    -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, 
    -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, 
    -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, 
    -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, 
    -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, 
    -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, 
    -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, 
    -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, 
    -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, 
    -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, 
    -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, 
    -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, 
    -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, 
    -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, 
    -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, 
    -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, -4.870118, 
    -4.870118, -4.870118,
  -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, 
    -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, 
    -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, 
    -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, 
    -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, 
    -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, 
    -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, 
    -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, 
    -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, 
    -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, 
    -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, 
    -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, 
    -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, 
    -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, 
    -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, 
    -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, 
    -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, 
    -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, 
    -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, 
    -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, 
    -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, 
    -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, 
    -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, 
    -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, 
    -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, 
    -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, 
    -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, 
    -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, 
    -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, 
    -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, -4.049516, 
    -4.049516, -4.049516,
  -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, 
    -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, 
    -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, 
    -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, 
    -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, 
    -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, 
    -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, 
    -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, 
    -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, 
    -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, 
    -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, 
    -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, 
    -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, 
    -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, 
    -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, 
    -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, 
    -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, 
    -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, 
    -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, 
    -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, 
    -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, 
    -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, 
    -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, 
    -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, 
    -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, 
    -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, 
    -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, 
    -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, 
    -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, 
    -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, -3.321665, 
    -3.321665, -3.321665,
  -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, 
    -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, 
    -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, 
    -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, 
    -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, 
    -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, 
    -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, 
    -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, 
    -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, 
    -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, 
    -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, 
    -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, 
    -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, 
    -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, 
    -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, 
    -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, 
    -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, 
    -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, 
    -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, 
    -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, 
    -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, 
    -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, 
    -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, 
    -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, 
    -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, 
    -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, 
    -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, 
    -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, 
    -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, 
    -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, -2.670094, 
    -2.670094, -2.670094,
  -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, 
    -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, 
    -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, 
    -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, 
    -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, 
    -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, 
    -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, 
    -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, 
    -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, 
    -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, 
    -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, 
    -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, 
    -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, 
    -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, 
    -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, 
    -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, 
    -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, 
    -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, 
    -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, 
    -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, 
    -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, 
    -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, 
    -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, 
    -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, 
    -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, 
    -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, 
    -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, 
    -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, 
    -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, 
    -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, -2.077874, 
    -2.077874, -2.077874,
  -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, 
    -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, 
    -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, 
    -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, 
    -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, 
    -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, 
    -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, 
    -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, 
    -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, 
    -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, 
    -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, 
    -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, 
    -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, 
    -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, 
    -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, 
    -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, 
    -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, 
    -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, 
    -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, 
    -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, 
    -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, 
    -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, 
    -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, 
    -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, 
    -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, 
    -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, 
    -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, 
    -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, 
    -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, 
    -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, -1.528546, 
    -1.528546, -1.528546,
  -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, 
    -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, 
    -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, 
    -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, 
    -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, 
    -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, 
    -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, 
    -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, 
    -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, 
    -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, 
    -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, 
    -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, 
    -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, 
    -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, 
    -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, 
    -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, 
    -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, 
    -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, 
    -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, 
    -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, 
    -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, 
    -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, 
    -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, 
    -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, 
    -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, 
    -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, 
    -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, 
    -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, 
    -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, 
    -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, -1.007058, 
    -1.007058, -1.007058,
  -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, 
    -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, 
    -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, 
    -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, 
    -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, 
    -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, 
    -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, 
    -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, 
    -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, 
    -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, 
    -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, 
    -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, 
    -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, 
    -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, 
    -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, 
    -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, 
    -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, 
    -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, 
    -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, 
    -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, 
    -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, 
    -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, 
    -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, 
    -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, 
    -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, 
    -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, 
    -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, 
    -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, 
    -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, 
    -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, -0.5006917, 
    -0.5006917, -0.5006917,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 
    0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 
    0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 
    0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 
    0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 
    0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 
    0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 
    0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 
    0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 
    0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 
    0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 
    0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 
    0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 
    0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 
    0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 
    0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 
    0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 
    0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 
    0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 
    0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 
    0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 
    0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 
    0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 
    0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 
    0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 
    0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 
    0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 
    0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 
    0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 
    0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 0.5006917, 
    0.5006917, 0.5006917,
  1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 
    1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 
    1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 
    1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 
    1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 
    1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 
    1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 
    1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 
    1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 
    1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 
    1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 
    1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 
    1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 
    1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 
    1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 
    1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 
    1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 
    1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 
    1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 
    1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 
    1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 
    1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 
    1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 
    1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 
    1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 
    1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058, 1.007058,
  1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 
    1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 
    1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 
    1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 
    1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 
    1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 
    1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 
    1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 
    1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 
    1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 
    1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 
    1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 
    1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 
    1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 
    1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 
    1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 
    1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 
    1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 
    1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 
    1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 
    1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 
    1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 
    1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 
    1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 
    1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 
    1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546, 1.528546,
  2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 
    2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 
    2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 
    2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 
    2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 
    2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 
    2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 
    2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 
    2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 
    2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 
    2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 
    2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 
    2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 
    2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 
    2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 
    2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 
    2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 
    2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 
    2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 
    2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 
    2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 
    2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 
    2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 
    2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 
    2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 
    2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874, 2.077874,
  2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 
    2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 
    2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 
    2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 
    2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 
    2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 
    2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 
    2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 
    2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 
    2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 
    2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 
    2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 
    2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 
    2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 
    2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 
    2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 
    2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 
    2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 
    2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 
    2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 
    2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 
    2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 
    2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 
    2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 
    2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 
    2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094, 2.670094,
  3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 
    3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 
    3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 
    3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 
    3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 
    3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 
    3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 
    3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 
    3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 
    3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 
    3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 
    3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 
    3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 
    3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 
    3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 
    3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 
    3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 
    3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 
    3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 
    3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 
    3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 
    3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 
    3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 
    3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 
    3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 
    3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665, 3.321665,
  4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 
    4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 
    4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 
    4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 
    4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 
    4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 
    4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 
    4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 
    4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 
    4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 
    4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 
    4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 
    4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 
    4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 
    4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 
    4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 
    4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 
    4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 
    4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 
    4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 
    4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 
    4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 
    4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 
    4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 
    4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 
    4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516, 4.049516,
  4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 
    4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 
    4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 
    4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 
    4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 
    4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 
    4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 
    4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 
    4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 
    4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 
    4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 
    4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 
    4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 
    4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 
    4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 
    4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 
    4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 
    4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 
    4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 
    4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 
    4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 
    4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 
    4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 
    4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 
    4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 
    4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118, 4.870118,
  5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 
    5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 
    5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 
    5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 
    5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 
    5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 
    5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 
    5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 
    5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 
    5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 
    5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 
    5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 
    5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 
    5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 
    5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 
    5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 
    5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 
    5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 
    5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 
    5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 
    5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 
    5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 
    5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 
    5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 
    5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 
    5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548, 5.798548,
  6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 
    6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 
    6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 
    6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 
    6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 
    6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 
    6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 
    6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 
    6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 
    6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 
    6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 
    6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 
    6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 
    6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 
    6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 
    6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 
    6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 
    6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 
    6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 
    6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 
    6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 
    6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 
    6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 
    6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 
    6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 
    6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561, 6.847561,
  8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 
    8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 
    8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 
    8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 
    8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 
    8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 
    8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 
    8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 
    8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 
    8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 
    8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 
    8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 
    8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 
    8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 
    8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 
    8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 
    8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 
    8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 
    8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 
    8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 
    8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 
    8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 
    8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 
    8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 
    8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 
    8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655, 8.026655,
  9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 
    9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 
    9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 
    9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 
    9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 
    9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 
    9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 
    9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 
    9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 
    9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 
    9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 
    9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 
    9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 
    9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 
    9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 
    9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 
    9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 
    9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 
    9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 
    9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 
    9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 
    9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 
    9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 
    9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 
    9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 
    9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137, 9.341137,
  10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 
    10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 
    10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 
    10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 
    10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 
    10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 
    10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 
    10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 
    10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 
    10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 
    10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 
    10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 
    10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 
    10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 
    10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 
    10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 
    10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 
    10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 
    10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 
    10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 
    10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 
    10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 
    10.7912, 10.7912, 10.7912, 10.7912, 10.7912, 10.7912,
  12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 
    12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 
    12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 
    12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 
    12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 
    12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 
    12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 
    12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 
    12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 
    12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 
    12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 
    12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 
    12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 
    12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 
    12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 
    12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 
    12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 
    12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 
    12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 
    12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 
    12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 
    12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 
    12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 
    12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 
    12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 
    12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097, 12.37097,
  14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 
    14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 
    14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 
    14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 
    14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 
    14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 
    14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 
    14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 
    14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 
    14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 
    14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 
    14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 
    14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 
    14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 
    14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 
    14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 
    14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 
    14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 
    14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 
    14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 
    14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 
    14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 
    14.0676, 14.0676, 14.0676, 14.0676, 14.0676, 14.0676,
  15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 
    15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 
    15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 
    15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 
    15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 
    15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 
    15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 
    15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 
    15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 
    15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 
    15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 
    15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 
    15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 
    15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 
    15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 
    15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 
    15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 
    15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 
    15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 
    15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 
    15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 
    15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 
    15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 
    15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 
    15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 
    15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032, 15.86032,
  17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 
    17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 
    17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 
    17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 
    17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 
    17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 
    17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 
    17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 
    17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 
    17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 
    17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 
    17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 
    17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 
    17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 
    17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 
    17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 
    17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 
    17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 
    17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 
    17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 
    17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 
    17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 
    17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 
    17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 
    17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 
    17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952, 17.71952,
  19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 
    19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 
    19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 
    19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 
    19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 
    19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 
    19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 
    19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 
    19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 
    19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 
    19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 
    19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 
    19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 
    19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 
    19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 
    19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 
    19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 
    19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 
    19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 
    19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 
    19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 
    19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 
    19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 
    19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 
    19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 
    19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579, 19.60579,
  21.47845, 21.47845, 21.47845, 21.47845, 21.47845, 21.47845, 21.47845, 
    21.47845, 21.47845, 21.47845, 21.47845, 21.47845, 21.47845, 21.47846, 
    21.47846, 21.47846, 21.47846, 21.47846, 21.47847, 21.47847, 21.47847, 
    21.47847, 21.47847, 21.47848, 21.47848, 21.47848, 21.47848, 21.47849, 
    21.47849, 21.47849, 21.47849, 21.47849, 21.4785, 21.4785, 21.4785, 
    21.4785, 21.4785, 21.47851, 21.47851, 21.47851, 21.47851, 21.47851, 
    21.47851, 21.47852, 21.47852, 21.47852, 21.47852, 21.47852, 21.47852, 
    21.47852, 21.47852, 21.47852, 21.47852, 21.47852, 21.47852, 21.47852, 
    21.47852, 21.47852, 21.47852, 21.47852, 21.47852, 21.47852, 21.47852, 
    21.47852, 21.47852, 21.47852, 21.47852, 21.47851, 21.47851, 21.47851, 
    21.47851, 21.47851, 21.47851, 21.47851, 21.47851, 21.47851, 21.4785, 
    21.4785, 21.4785, 21.4785, 21.4785, 21.4785, 21.4785, 21.4785, 21.4785, 
    21.4785, 21.4785, 21.4785, 21.4785, 21.4785, 21.4785, 21.4785, 21.4785, 
    21.4785, 21.4785, 21.4785, 21.4785, 21.4785, 21.4785, 21.4785, 21.4785, 
    21.4785, 21.4785, 21.4785, 21.4785, 21.4785, 21.4785, 21.47851, 21.47851, 
    21.47851, 21.47851, 21.47851, 21.47851, 21.47851, 21.47851, 21.47851, 
    21.47852, 21.47852, 21.47852, 21.47852, 21.47852, 21.47852, 21.47852, 
    21.47852, 21.47852, 21.47852, 21.47852, 21.47852, 21.47852, 21.47852, 
    21.47852, 21.47852, 21.47852, 21.47852, 21.47852, 21.47852, 21.47852, 
    21.47852, 21.47852, 21.47846, 21.47846, 21.47846, 21.47846, 21.47846, 
    21.47846, 21.47846, 21.47846, 21.47846, 21.47846, 21.47846, 21.47846, 
    21.47846, 21.47846, 21.47846, 21.47846, 21.47846, 21.47846, 21.47846, 
    21.47846, 21.47846, 21.47846, 21.47846, 21.47846, 21.47846, 21.47846, 
    21.47846, 21.47846, 21.47846, 21.47846, 21.47846, 21.47845, 21.47845, 
    21.47845, 21.47845, 21.47845, 21.47845, 21.47845, 21.47845, 21.47845, 
    21.47845, 21.47845, 21.47845,
  23.32185, 23.32184, 23.32185, 23.32186, 23.32189, 23.32193, 23.32198, 
    23.32204, 23.32212, 23.3222, 23.32229, 23.3224, 23.32251, 23.32263, 
    23.32276, 23.32289, 23.32304, 23.32319, 23.32334, 23.3235, 23.32367, 
    23.32384, 23.32401, 23.32419, 23.32437, 23.32455, 23.32473, 23.32491, 
    23.32509, 23.32527, 23.32545, 23.32562, 23.32579, 23.32596, 23.32612, 
    23.32628, 23.32643, 23.32658, 23.32672, 23.32685, 23.32697, 23.32709, 
    23.3272, 23.3273, 23.32739, 23.32747, 23.32755, 23.32761, 23.32767, 
    23.32772, 23.32775, 23.32778, 23.3278, 23.32781, 23.32782, 23.32781, 
    23.3278, 23.32778, 23.32775, 23.32771, 23.32767, 23.32762, 23.32756, 
    23.32751, 23.32744, 23.32737, 23.3273, 23.32722, 23.32714, 23.32706, 
    23.32698, 23.3269, 23.32682, 23.32673, 23.32665, 23.32657, 23.32649, 
    23.32642, 23.32635, 23.32627, 23.32621, 23.32615, 23.32609, 23.32604, 
    23.32599, 23.32595, 23.32591, 23.32589, 23.32586, 23.32585, 23.32584, 
    23.32583, 23.32584, 23.32585, 23.32586, 23.32589, 23.32591, 23.32595, 
    23.32599, 23.32604, 23.32609, 23.32615, 23.32621, 23.32627, 23.32635, 
    23.32642, 23.32649, 23.32657, 23.32665, 23.32673, 23.32682, 23.3269, 
    23.32698, 23.32706, 23.32714, 23.32722, 23.3273, 23.32737, 23.32744, 
    23.32751, 23.32756, 23.32762, 23.32767, 23.32771, 23.32775, 23.32778, 
    23.3278, 23.32781, 23.32782, 23.32781, 23.3278, 23.32778, 23.32775, 
    23.32772, 23.32767, 23.32761, 23.32755, 23.32747, 23.32739, 23.32289, 
    23.32289, 23.32289, 23.32289, 23.32289, 23.32289, 23.32289, 23.32289, 
    23.32289, 23.32289, 23.32289, 23.32289, 23.32289, 23.32289, 23.32289, 
    23.32289, 23.32289, 23.32289, 23.32289, 23.32289, 23.32289, 23.32289, 
    23.32289, 23.32289, 23.32289, 23.32289, 23.32289, 23.32289, 23.32289, 
    23.32276, 23.32263, 23.32251, 23.3224, 23.32229, 23.3222, 23.32212, 
    23.32204, 23.32198, 23.32193, 23.32189, 23.32186, 23.32185, 23.32184,
  25.12383, 25.1238, 25.12383, 25.12391, 25.12405, 25.12425, 25.12449, 
    25.12479, 25.12514, 25.12555, 25.126, 25.12649, 25.12704, 25.12762, 
    25.12824, 25.1289, 25.1296, 25.13033, 25.13109, 25.13187, 25.13268, 
    25.1335, 25.13435, 25.1352, 25.13607, 25.13694, 25.13782, 25.1387, 
    25.13957, 25.14044, 25.14129, 25.14214, 25.14297, 25.14377, 25.14456, 
    25.14532, 25.14606, 25.14676, 25.14744, 25.14808, 25.14868, 25.14925, 
    25.14978, 25.15026, 25.15071, 25.15111, 25.15147, 25.15178, 25.15206, 
    25.15228, 25.15247, 25.15261, 25.1527, 25.15276, 25.15277, 25.15274, 
    25.15267, 25.15257, 25.15243, 25.15225, 25.15204, 25.15181, 25.15154, 
    25.15125, 25.15094, 25.1506, 25.15025, 25.14989, 25.14951, 25.14912, 
    25.14872, 25.14832, 25.14792, 25.14752, 25.14712, 25.14673, 25.14635, 
    25.14598, 25.14563, 25.14529, 25.14497, 25.14467, 25.14439, 25.14414, 
    25.14391, 25.14371, 25.14354, 25.1434, 25.14329, 25.14321, 25.14316, 
    25.14315, 25.14316, 25.14321, 25.14329, 25.1434, 25.14354, 25.14371, 
    25.14391, 25.14414, 25.14439, 25.14467, 25.14497, 25.14529, 25.14563, 
    25.14598, 25.14635, 25.14673, 25.14712, 25.14752, 25.14792, 25.14832, 
    25.14872, 25.14912, 25.14951, 25.14989, 25.15025, 25.1506, 25.15094, 
    25.15125, 25.15154, 25.15181, 25.15204, 25.15225, 25.15243, 25.15257, 
    25.15267, 25.15274, 25.15277, 25.15276, 25.1527, 25.15261, 25.15247, 
    25.15228, 25.15206, 25.15178, 25.15147, 25.15111, 25.15071, 25.1289, 
    25.1289, 25.1289, 25.1289, 25.1289, 25.1289, 25.1289, 25.1289, 25.1289, 
    25.1289, 25.1289, 25.1289, 25.1289, 25.1289, 29.51136, 29.51136, 
    29.51136, 29.51136, 29.51136, 29.51136, 29.51136, 29.51136, 29.51136, 
    29.51136, 29.51136, 29.51136, 29.51136, 29.51136, 29.51136, 29.51136, 
    29.51136, 25.1238, 25.1238, 25.1238, 25.1238, 25.1238, 25.1238, 25.1238, 
    29.51136, 29.51136, 29.51136, 29.51136, 25.1238,
  26.87389, 26.87381, 26.87389, 26.87411, 26.87449, 26.87502, 26.87569, 
    26.8765, 26.87746, 26.87856, 26.87978, 26.88113, 26.88261, 26.8842, 
    26.88589, 26.8877, 26.88959, 26.89157, 26.89363, 26.89577, 26.89796, 
    26.90021, 26.90251, 26.90484, 26.9072, 26.90957, 26.91196, 26.91434, 
    26.91672, 26.91907, 26.9214, 26.92369, 26.92595, 26.92814, 26.93028, 
    26.93235, 26.93435, 26.93627, 26.9381, 26.93984, 26.94148, 26.94302, 
    26.94445, 26.94577, 26.94698, 26.94807, 26.94905, 26.9499, 26.95064, 
    26.95126, 26.95175, 26.95213, 26.95239, 26.95253, 26.95256, 26.95248, 
    26.9523, 26.95201, 26.95163, 26.95115, 26.95058, 26.94993, 26.94921, 
    26.94842, 26.94757, 26.94666, 26.9457, 26.9447, 26.94366, 26.9426, 
    26.94152, 26.94043, 26.93934, 26.93825, 26.93717, 26.93611, 26.93507, 
    26.93406, 26.9331, 26.93217, 26.9313, 26.93049, 26.92974, 26.92905, 
    26.92843, 26.92789, 26.92742, 26.92704, 26.92673, 26.92652, 26.92639, 
    26.92634, 26.92639, 26.92652, 26.92673, 26.92704, 26.92742, 26.92789, 
    26.92843, 26.92905, 26.92974, 26.93049, 26.9313, 26.93217, 26.9331, 
    26.93406, 26.93507, 26.93611, 26.93717, 26.93825, 26.93934, 26.94043, 
    26.94152, 26.9426, 26.94366, 26.9447, 26.9457, 26.94666, 26.94757, 
    26.94842, 26.94921, 26.94993, 26.95058, 26.95115, 26.95163, 26.95201, 
    26.9523, 26.95248, 26.95256, 26.95253, 26.95239, 26.95213, 26.95175, 
    26.95126, 26.95064, 26.9499, 26.94905, 26.94807, 26.94698, 26.8877, 
    26.8877, 26.8877, 26.8877, 26.8877, 26.8877, 26.8877, 26.8877, 26.8877, 
    26.8877, 26.8877, 26.8877, 26.8877, 26.8877, 30.51136, 30.51136, 
    30.51136, 30.51136, 30.51136, 30.51136, 30.51136, 30.51136, 30.51136, 
    30.51136, 30.51136, 30.51136, 30.51136, 30.51136, 30.51136, 30.51136, 
    30.51136, 30.51136, 30.51136, 30.51136, 30.51136, 30.51136, 30.51136, 
    30.51136, 30.51136, 30.51136, 30.51136, 30.51136, 26.87381,
  28.56264, 28.56248, 28.56264, 28.56311, 28.5639, 28.56499, 28.5664, 
    28.5681, 28.5701, 28.57238, 28.57494, 28.57776, 28.58083, 28.58415, 
    28.58769, 28.59145, 28.5954, 28.59954, 28.60384, 28.60829, 28.61286, 
    28.61755, 28.62234, 28.6272, 28.63211, 28.63706, 28.64203, 28.647, 
    28.65194, 28.65685, 28.6617, 28.66648, 28.67117, 28.67574, 28.68019, 
    28.68451, 28.68867, 28.69266, 28.69646, 28.70008, 28.7035, 28.7067, 
    28.70967, 28.71242, 28.71493, 28.7172, 28.71923, 28.72101, 28.72253, 
    28.72381, 28.72484, 28.72562, 28.72615, 28.72645, 28.72651, 28.72634, 
    28.72595, 28.72534, 28.72453, 28.72353, 28.72235, 28.721, 28.71949, 
    28.71783, 28.71605, 28.71415, 28.71215, 28.71006, 28.7079, 28.70569, 
    28.70343, 28.70116, 28.69887, 28.69659, 28.69434, 28.69212, 28.68996, 
    28.68786, 28.68584, 28.68391, 28.68209, 28.68039, 28.67882, 28.67738, 
    28.67609, 28.67496, 28.67399, 28.67318, 28.67255, 28.6721, 28.67183, 
    28.67173, 28.67183, 28.6721, 28.67255, 28.67318, 28.67399, 28.67496, 
    28.67609, 28.67738, 28.67882, 28.68039, 28.68209, 28.68391, 28.68584, 
    28.68786, 28.68996, 28.69212, 28.69434, 28.69659, 28.69887, 28.70116, 
    28.70343, 28.70569, 28.7079, 28.71006, 28.71215, 28.71415, 28.71605, 
    28.71783, 28.71949, 28.721, 28.72235, 28.72353, 28.72453, 28.72534, 
    28.72595, 28.72634, 28.72651, 28.72645, 28.72615, 28.72562, 28.72484, 
    28.72381, 28.72253, 28.72101, 28.71923, 28.7172, 28.71493, 28.59145, 
    28.59145, 28.59145, 28.59145, 28.59145, 28.59145, 28.59145, 28.59145, 
    28.59145, 28.59145, 31.51136, 31.51136, 31.51136, 31.51136, 31.51136, 
    31.51136, 31.51136, 31.51136, 31.51136, 31.51136, 31.51136, 31.51136, 
    31.51136, 31.51136, 31.51136, 31.51136, 31.51136, 31.51136, 31.51136, 
    31.51136, 31.51136, 31.51136, 31.51136, 31.51136, 31.51136, 31.51136, 
    31.51136, 31.51136, 31.51136, 31.51136, 31.51136, 31.51136, 28.56248,
  30.18224, 30.18196, 30.18224, 30.18308, 30.18449, 30.18645, 30.18896, 
    30.192, 30.19556, 30.19963, 30.2042, 30.20924, 30.21473, 30.22064, 
    30.22697, 30.23367, 30.24072, 30.2481, 30.25577, 30.2637, 30.27187, 
    30.28023, 30.28876, 30.29741, 30.30617, 30.31499, 30.32384, 30.33269, 
    30.3415, 30.35024, 30.35888, 30.36738, 30.37572, 30.38386, 30.39178, 
    30.39945, 30.40685, 30.41394, 30.42071, 30.42714, 30.4332, 30.43889, 
    30.44418, 30.44906, 30.45352, 30.45755, 30.46114, 30.46429, 30.467, 
    30.46926, 30.47108, 30.47246, 30.4734, 30.47391, 30.47401, 30.47369, 
    30.47299, 30.4719, 30.47046, 30.46867, 30.46655, 30.46413, 30.46144, 
    30.45848, 30.45529, 30.4519, 30.44833, 30.4446, 30.44075, 30.43679, 
    30.43277, 30.42871, 30.42463, 30.42056, 30.41654, 30.41258, 30.40871, 
    30.40497, 30.40136, 30.39792, 30.39468, 30.39164, 30.38882, 30.38626, 
    30.38396, 30.38193, 30.38019, 30.37876, 30.37763, 30.37682, 30.37633, 
    30.37617, 30.37633, 30.37682, 30.37763, 30.37876, 30.38019, 30.38193, 
    30.38396, 30.38626, 30.38882, 30.39164, 30.39468, 30.39792, 30.40136, 
    30.40497, 30.40871, 30.41258, 30.41654, 30.42056, 30.42463, 30.42871, 
    30.43277, 30.43679, 30.44075, 30.4446, 30.44833, 30.4519, 30.45529, 
    30.45848, 30.46144, 30.46413, 30.46655, 30.46867, 30.47046, 30.4719, 
    30.47299, 30.47369, 30.47401, 30.47391, 30.4734, 30.47246, 30.47108, 
    30.46926, 30.467, 30.46429, 30.46114, 30.45755, 30.45352, 30.4235, 
    32.51136, 32.51136, 32.51136, 32.51136, 32.51136, 32.51136, 32.51136, 
    32.51136, 32.51136, 32.51136, 32.51136, 32.51136, 32.51136, 32.51136, 
    32.51136, 32.51136, 32.51136, 32.51136, 32.51136, 32.51136, 32.51136, 
    32.51136, 32.51136, 32.51136, 32.51136, 32.51136, 32.51136, 32.51136, 
    32.51136, 32.51136, 32.51136, 32.51136, 32.51136, 32.51136, 32.51136, 
    32.51136, 32.51136, 32.51136, 32.51136, 32.51136, 32.51136, 30.18196,
  31.7265, 31.7265, 31.7265, 31.72786, 31.73012, 31.73328, 31.73732, 
    31.74221, 31.74796, 31.75451, 31.76186, 31.76997, 31.7788, 31.78833, 
    31.7985, 31.80928, 31.82063, 31.83249, 31.84483, 31.85758, 31.8707, 
    31.88414, 31.89784, 31.91175, 31.92581, 31.93997, 31.95418, 31.96838, 
    31.98251, 31.99653, 32.01038, 32.02401, 32.03738, 32.05043, 32.06312, 
    32.07541, 32.08725, 32.09861, 32.10945, 32.11974, 32.12944, 32.13854, 
    32.147, 32.1548, 32.16193, 32.16837, 32.17411, 32.17914, 32.18345, 
    32.18706, 32.18995, 32.19213, 32.19363, 32.19443, 32.19456, 32.19404, 
    32.19289, 32.19113, 32.1888, 32.18591, 32.1825, 32.1786, 32.17426, 
    32.16951, 32.16438, 32.15892, 32.15317, 32.14717, 32.14097, 32.13462, 
    32.12815, 32.12161, 32.11505, 32.10851, 32.10203, 32.09566, 32.08944, 
    32.08341, 32.07761, 32.07208, 32.06685, 32.06195, 32.05743, 32.0533, 
    32.04959, 32.04633, 32.04353, 32.04122, 32.03941, 32.0381, 32.03732, 
    32.03705, 32.03732, 32.0381, 32.03941, 32.04122, 32.04353, 32.04633, 
    32.04959, 32.0533, 32.05743, 32.06195, 32.06685, 32.07208, 32.07761, 
    32.08341, 32.08944, 32.09566, 32.10203, 32.10851, 32.11505, 32.12161, 
    32.12815, 32.13462, 32.14097, 32.14717, 32.15317, 32.15892, 32.16438, 
    32.16951, 32.17426, 32.1786, 32.1825, 32.18591, 32.1888, 32.19113, 
    32.19289, 32.19404, 32.19456, 32.19443, 32.19363, 32.19213, 32.18995, 
    32.18706, 32.18345, 32.17914, 32.17411, 32.29265, 32.49802, 32.60139, 
    33.51136, 33.51136, 33.51136, 33.51136, 33.51136, 33.51136, 33.51136, 
    33.51136, 33.51136, 33.51136, 33.51136, 33.51136, 33.51136, 33.51136, 
    33.51136, 33.51136, 33.51136, 33.51136, 33.51136, 33.51136, 33.51136, 
    33.51136, 33.51136, 33.51136, 33.51136, 33.51136, 33.51136, 33.51136, 
    33.51136, 33.51136, 33.51136, 33.51136, 33.51136, 33.51136, 33.51136, 
    33.51136, 33.51136, 33.51136, 33.51136, 33.51136, 33.51136, 33.51136,
  33.19087, 33.19087, 33.19087, 33.19291, 33.1963, 33.20102, 33.20706, 
    33.21439, 33.22298, 33.23279, 33.24378, 33.2559, 33.26911, 33.28334, 
    33.29855, 33.31466, 33.33161, 33.34933, 33.36774, 33.38678, 33.40636, 
    33.42641, 33.44684, 33.46758, 33.48855, 33.50965, 33.53082, 33.55197, 
    33.57301, 33.59388, 33.61449, 33.63478, 33.65466, 33.67406, 33.69292, 
    33.71119, 33.72878, 33.74565, 33.76175, 33.77702, 33.79142, 33.80491, 
    33.81745, 33.82902, 33.83958, 33.84912, 33.85762, 33.86506, 33.87144, 
    33.87677, 33.88103, 33.88425, 33.88643, 33.88759, 33.88775, 33.88695, 
    33.8852, 33.88256, 33.87906, 33.87473, 33.86963, 33.86381, 33.85732, 
    33.85021, 33.84256, 33.8344, 33.82582, 33.81686, 33.80761, 33.79812, 
    33.78846, 33.77869, 33.76889, 33.75912, 33.74945, 33.73994, 33.73064, 
    33.72164, 33.71297, 33.7047, 33.69689, 33.68958, 33.68281, 33.67663, 
    33.67109, 33.66621, 33.66203, 33.65857, 33.65586, 33.65392, 33.65274, 
    33.65235, 33.65274, 33.65392, 33.65586, 33.65857, 33.66203, 33.66621, 
    33.67109, 33.67663, 33.68281, 33.68958, 33.69689, 33.7047, 33.71297, 
    33.72164, 33.73064, 33.73994, 33.74945, 33.75912, 33.76889, 33.77869, 
    33.78846, 33.79812, 33.80761, 33.81686, 33.82582, 33.8344, 33.84256, 
    33.85021, 33.85732, 33.86381, 33.86963, 33.87473, 33.87906, 33.88256, 
    33.8852, 33.88695, 33.88775, 33.88759, 33.88643, 33.88425, 33.88103, 
    33.87677, 33.87144, 33.86506, 33.85762, 34.1845, 34.4024, 34.51136, 
    34.51136, 34.51136, 34.51136, 34.51136, 34.51136, 34.51136, 34.51136, 
    34.51136, 34.51136, 34.51136, 34.51136, 34.51136, 34.51136, 34.51136, 
    34.51136, 34.51136, 34.51136, 34.51136, 34.51136, 34.51136, 34.51136, 
    34.51136, 34.51136, 34.51136, 34.51136, 34.51136, 34.51136, 34.51136, 
    34.51136, 34.51136, 34.51136, 34.51136, 34.51136, 34.51136, 34.51136, 
    34.51136, 34.51136, 34.51136, 34.51136, 34.51136, 34.51136, 34.51136,
  34.57241, 34.57241, 34.57241, 34.5753, 34.5801, 34.58679, 34.59534, 
    34.60572, 34.61788, 34.63176, 34.64732, 34.66447, 34.68316, 34.70329, 
    34.72479, 34.74757, 34.77152, 34.79655, 34.82256, 34.84944, 34.87708, 
    34.90536, 34.93419, 34.96343, 34.99298, 35.02272, 35.05253, 35.0823, 
    35.11193, 35.14129, 35.17028, 35.1988, 35.22674, 35.25401, 35.2805, 
    35.30614, 35.33084, 35.35451, 35.37709, 35.3985, 35.41869, 35.43759, 
    35.45516, 35.47136, 35.48614, 35.49948, 35.51136, 35.52176, 35.53067, 
    35.53809, 35.54403, 35.54848, 35.55149, 35.55307, 35.55325, 35.55207, 
    35.54957, 35.5458, 35.54083, 35.5347, 35.52749, 35.51926, 35.51009, 
    35.50006, 35.48924, 35.47773, 35.46561, 35.45298, 35.43991, 35.42651, 
    35.41288, 35.39909, 35.38526, 35.37146, 35.3578, 35.34436, 35.33124, 
    35.31851, 35.30627, 35.29458, 35.28354, 35.27319, 35.26363, 35.2549, 
    35.24706, 35.24016, 35.23425, 35.22936, 35.22552, 35.22277, 35.22111, 
    35.22055, 35.22111, 35.22277, 35.22552, 35.22936, 35.23425, 35.24016, 
    35.24706, 35.2549, 35.26363, 35.27319, 35.28354, 35.29458, 35.30627, 
    35.31851, 35.33124, 35.34436, 35.3578, 35.37146, 35.38526, 35.39909, 
    35.41288, 35.42651, 35.43991, 35.45298, 35.46561, 35.47773, 35.48924, 
    35.50006, 35.51009, 35.51926, 35.52749, 35.5347, 35.54083, 35.5458, 
    35.54957, 35.55207, 35.55325, 35.55307, 35.55149, 35.54848, 35.54403, 
    35.53809, 35.53067, 35.52176, 35.51136, 35.51136, 35.51136, 35.51136, 
    35.51136, 35.51136, 35.51136, 35.51136, 35.51136, 35.51136, 35.51136, 
    35.51136, 35.51136, 35.51136, 35.51136, 35.51136, 35.51136, 35.51136, 
    35.51136, 35.51136, 35.51136, 35.51136, 35.51136, 35.51136, 35.51136, 
    35.51136, 35.51136, 35.51136, 35.51136, 35.51136, 35.51136, 35.51136, 
    35.51136, 35.51136, 35.51136, 35.51136, 35.51136, 35.51136, 35.51136, 
    35.51136, 35.51136, 35.51136, 35.51136, 35.51136, 35.51136, 35.51136,
  35.86965, 35.86965, 35.86965, 35.87357, 35.88008, 35.88916, 35.90077, 
    35.91485, 35.93134, 35.95018, 35.97127, 35.99452, 36.01984, 36.04712, 
    36.07624, 36.10707, 36.1395, 36.17336, 36.20854, 36.24488, 36.28223, 
    36.32044, 36.35936, 36.39883, 36.43869, 36.47879, 36.51899, 36.5591, 
    36.599, 36.63853, 36.67755, 36.71591, 36.75348, 36.79013, 36.82573, 
    36.86016, 36.89332, 36.92509, 36.95538, 36.98409, 37.01115, 37.03647, 
    37.06001, 37.08168, 37.10147, 37.11931, 37.13518, 37.14907, 37.16095, 
    37.17084, 37.17873, 37.18464, 37.1886, 37.19064, 37.1908, 37.18914, 
    37.1857, 37.18057, 37.17381, 37.1655, 37.15573, 37.1446, 37.13219, 
    37.11863, 37.10402, 37.08847, 37.0721, 37.05502, 37.03738, 37.01927, 
    37.00085, 36.98222, 36.96352, 36.94487, 36.9264, 36.90823, 36.89049, 
    36.87327, 36.85671, 36.8409, 36.82595, 36.81196, 36.79901, 36.78719, 
    36.77658, 36.76724, 36.75924, 36.75261, 36.74742, 36.74369, 36.74144, 
    36.74068, 36.74144, 36.74369, 36.74742, 36.75261, 36.75924, 36.76724, 
    36.77658, 36.78719, 36.79901, 36.81196, 36.82595, 36.8409, 36.85671, 
    36.87327, 36.89049, 36.90823, 36.9264, 36.94487, 36.96352, 36.98222, 
    37.00085, 37.01927, 37.03738, 37.05502, 37.0721, 37.08847, 37.10402, 
    37.11863, 37.13219, 37.1446, 37.15573, 37.1655, 37.17381, 37.18057, 
    37.1857, 37.18914, 37.1908, 37.19064, 37.1886, 37.18464, 37.17873, 
    37.17084, 37.16095, 37.14907, 37.13518, 36.8233, 36.6153, 36.51136, 
    36.51136, 36.51136, 36.51136, 36.51136, 36.51136, 36.51136, 36.51136, 
    36.51136, 36.51136, 36.51136, 36.51136, 36.51136, 36.51136, 36.51136, 
    36.51136, 36.51136, 36.51136, 36.51136, 36.51136, 36.51136, 36.51136, 
    36.51136, 36.51136, 36.51136, 36.51136, 36.51136, 36.51136, 36.51136, 
    36.51136, 36.51136, 36.51136, 36.51136, 36.51136, 36.51136, 36.51136, 
    36.51136, 36.51136, 36.51136, 36.51136, 36.51136, 36.51136, 36.51136,
  37.08244, 37.08244, 37.08244, 37.08759, 37.09613, 37.10804, 37.12326, 
    37.14173, 37.16335, 37.18803, 37.21567, 37.24614, 37.2793, 37.31501, 
    37.35311, 37.39344, 37.43583, 37.48009, 37.52604, 37.57349, 37.62224, 
    37.67208, 37.72283, 37.77426, 37.82619, 37.8784, 37.9307, 37.98288, 
    38.03474, 38.08611, 38.13678, 38.18658, 38.23533, 38.28286, 38.32901, 
    38.37362, 38.41656, 38.45769, 38.49688, 38.53402, 38.569, 38.60173, 
    38.63213, 38.66012, 38.68564, 38.70865, 38.7291, 38.74697, 38.76226, 
    38.77495, 38.78506, 38.7926, 38.79762, 38.80014, 38.80024, 38.79797, 
    38.79341, 38.78664, 38.77777, 38.76689, 38.75411, 38.73957, 38.72338, 
    38.70568, 38.68661, 38.66633, 38.64498, 38.62271, 38.59969, 38.57608, 
    38.55204, 38.52774, 38.50335, 38.47901, 38.4549, 38.43119, 38.40801, 
    38.38553, 38.3639, 38.34324, 38.32371, 38.30542, 38.28849, 38.27304, 
    38.25917, 38.24695, 38.23648, 38.22782, 38.22103, 38.21614, 38.2132, 
    38.21221, 38.2132, 38.21614, 38.22103, 38.22782, 38.23648, 38.24695, 
    38.25917, 38.27304, 38.28849, 38.30542, 38.32371, 38.34324, 38.3639, 
    38.38553, 38.40801, 38.43119, 38.4549, 38.47901, 38.50335, 38.52774, 
    38.55204, 38.57608, 38.59969, 38.62271, 38.64498, 38.66633, 38.68661, 
    38.70568, 38.72338, 38.73957, 38.75411, 38.76689, 38.77777, 38.78664, 
    38.79341, 38.79797, 38.80024, 38.80014, 38.79762, 38.7926, 38.78506, 
    38.77495, 38.76226, 38.74697, 38.7291, 38.31762, 37.77465, 37.56333, 
    37.51136, 37.51136, 37.51136, 37.51136, 37.51136, 37.51136, 37.51136, 
    37.51136, 37.51136, 37.51136, 37.51136, 37.51136, 37.51136, 37.51136, 
    37.51136, 37.51136, 37.51136, 37.51136, 37.51136, 37.51136, 37.51136, 
    37.51136, 37.51136, 37.51136, 37.51136, 37.51136, 37.51136, 37.51136, 
    37.51136, 37.51136, 37.51136, 37.51136, 37.51136, 37.51136, 37.51136, 
    37.51136, 37.51136, 37.51136, 37.51136, 37.51136, 37.51136, 37.51136,
  38.21178, 38.20959, 38.21178, 38.21835, 38.22926, 38.24445, 38.26387, 
    38.28742, 38.31499, 38.34646, 38.38168, 38.42049, 38.46272, 38.50817, 
    38.55665, 38.60794, 38.66182, 38.71805, 38.7764, 38.83661, 38.89844, 
    38.96162, 39.02591, 39.09104, 39.15675, 39.22279, 39.28889, 39.35482, 
    39.42031, 39.48512, 39.54903, 39.61181, 39.67323, 39.73308, 39.79117, 
    39.8473, 39.90129, 39.95298, 40.00221, 40.04884, 40.09274, 40.13379, 
    40.1719, 40.20697, 40.23892, 40.26771, 40.29328, 40.31561, 40.33467, 
    40.35047, 40.36302, 40.37234, 40.37849, 40.38151, 40.38147, 40.37846, 
    40.37257, 40.3639, 40.35258, 40.33873, 40.3225, 40.30404, 40.2835, 
    40.26106, 40.2369, 40.21119, 40.18414, 40.15593, 40.12676, 40.09684, 
    40.06638, 40.03557, 40.00464, 39.97379, 39.94321, 39.91313, 39.88372, 
    39.8552, 39.82774, 39.80152, 39.77671, 39.75348, 39.73198, 39.71235, 
    39.69472, 39.6792, 39.66589, 39.65487, 39.64623, 39.64002, 39.63628, 
    39.63503, 39.63628, 39.64002, 39.64623, 39.65487, 39.66589, 39.6792, 
    39.69472, 39.71235, 39.73198, 39.75348, 39.77671, 39.80152, 39.82774, 
    39.8552, 39.88372, 39.91313, 39.94321, 39.97379, 40.00464, 40.03557, 
    40.06638, 40.09684, 40.12676, 40.15593, 40.18414, 40.21119, 40.2369, 
    40.26106, 40.2835, 40.30404, 40.3225, 40.33873, 40.35258, 40.3639, 
    40.37257, 40.37846, 40.38147, 40.38151, 40.37849, 40.37234, 40.36302, 
    40.35047, 40.33467, 40.31561, 40.29328, 40.02278, 39.67334, 39.53127, 
    38.51136, 38.51136, 38.51136, 38.51136, 38.51136, 38.51136, 38.51136, 
    38.51136, 38.51136, 38.51136, 38.51136, 38.51136, 38.51136, 38.51136, 
    38.51136, 38.51136, 38.51136, 38.51136, 38.51136, 38.51136, 38.51136, 
    38.51136, 38.51136, 38.51136, 38.51136, 38.51136, 38.51136, 38.51136, 
    38.51136, 38.51136, 38.51136, 38.51136, 38.51136, 38.51136, 38.51136, 
    38.51136, 38.51136, 38.51136, 38.51136, 38.51136, 38.51136, 38.20959,
  39.25962, 39.25689, 39.25962, 39.26781, 39.28142, 39.30037, 39.32459, 
    39.35395, 39.38831, 39.42751, 39.47137, 39.51969, 39.57223, 39.62875, 
    39.68901, 39.75273, 39.81962, 39.88939, 39.96174, 40.03636, 40.11293, 
    40.19114, 40.27065, 40.35115, 40.43233, 40.51385, 40.5954, 40.67668, 
    40.75737, 40.83719, 40.91585, 40.99306, 41.06856, 41.14209, 41.21342, 
    41.2823, 41.34853, 41.4119, 41.47222, 41.52932, 41.58306, 41.63328, 
    41.67986, 41.72271, 41.76173, 41.79684, 41.82801, 41.85519, 41.87837, 
    41.89754, 41.91273, 41.92396, 41.93128, 41.93477, 41.93451, 41.9306, 
    41.92316, 41.91231, 41.8982, 41.88099, 41.86085, 41.83797, 41.81253, 
    41.78476, 41.75486, 41.72306, 41.68959, 41.6547, 41.61862, 41.58162, 
    41.54393, 41.50581, 41.46753, 41.42934, 41.39149, 41.35423, 41.31781, 
    41.28247, 41.24844, 41.21594, 41.18518, 41.15638, 41.12971, 41.10535, 
    41.08347, 41.06421, 41.04768, 41.03401, 41.02329, 41.01558, 41.01093, 
    41.00937, 41.01093, 41.01558, 41.02329, 41.03401, 41.04768, 41.06421, 
    41.08347, 41.10535, 41.12971, 41.15638, 41.18518, 41.21594, 41.24844, 
    41.28247, 41.31781, 41.35423, 41.39149, 41.42934, 41.46753, 41.50581, 
    41.54393, 41.58162, 41.61862, 41.6547, 41.68959, 41.72306, 41.75486, 
    41.78476, 41.81253, 41.83797, 41.86085, 41.88099, 41.8982, 41.91231, 
    41.92316, 41.9306, 41.93451, 41.93477, 41.93128, 41.92396, 41.91273, 
    41.89754, 41.87837, 41.85519, 41.82801, 41.79684, 41.76173, 41.72271, 
    39.51136, 39.51136, 39.51136, 39.51136, 39.51136, 39.51136, 39.51136, 
    39.51136, 39.51136, 39.51136, 39.51136, 39.51136, 39.51136, 39.51136, 
    39.51136, 39.51136, 39.51136, 39.51136, 39.51136, 39.51136, 39.51136, 
    39.51136, 39.51136, 39.51136, 39.51136, 39.51136, 39.51136, 39.51136, 
    39.51136, 39.51136, 39.51136, 39.51136, 39.51136, 39.51136, 39.51136, 
    39.51136, 39.51136, 39.51136, 39.51136, 39.51136, 39.51136, 39.25689,
  40.22866, 40.22532, 40.22866, 40.23869, 40.25534, 40.27854, 40.30817, 
    40.34407, 40.38608, 40.43399, 40.48757, 40.54655, 40.61066, 40.67959, 
    40.75303, 40.83063, 40.91205, 40.99691, 41.08485, 41.17548, 41.26842, 
    41.36327, 41.45964, 41.55713, 41.65537, 41.75396, 41.85252, 41.95068, 
    42.04807, 42.14433, 42.23914, 42.33214, 42.42303, 42.51149, 42.59725, 
    42.68003, 42.75956, 42.83562, 42.90799, 42.97646, 43.04084, 43.10098, 
    43.15673, 43.20798, 43.25461, 43.29654, 43.33372, 43.3661, 43.39367, 
    43.41643, 43.43439, 43.44759, 43.45612, 43.46003, 43.45943, 43.45446, 
    43.44523, 43.43191, 43.41467, 43.3937, 43.36921, 43.34142, 43.31055, 
    43.27687, 43.24062, 43.20207, 43.16151, 43.11922, 43.0755, 43.03064, 
    42.98496, 42.93875, 42.89233, 42.84602, 42.8001, 42.75489, 42.71069, 
    42.66777, 42.62645, 42.58697, 42.5496, 42.51459, 42.48217, 42.45256, 
    42.42595, 42.40251, 42.38241, 42.36578, 42.35273, 42.34334, 42.33768, 
    42.33579, 42.33768, 42.34334, 42.35273, 42.36578, 42.38241, 42.40251, 
    42.42595, 42.45256, 42.48217, 42.51459, 42.5496, 42.58697, 42.62645, 
    42.66777, 42.71069, 42.75489, 42.8001, 42.84602, 42.89233, 42.93875, 
    42.98496, 43.03064, 43.0755, 43.11922, 43.16151, 43.20207, 43.24062, 
    43.27687, 43.31055, 43.34142, 43.36921, 43.3937, 43.41467, 43.43191, 
    43.44523, 43.45446, 43.45943, 43.46003, 43.45612, 43.44759, 43.43439, 
    43.41643, 43.39367, 43.3661, 43.33372, 43.29654, 43.25461, 43.20798, 
    43.15673, 43.10098, 43.20098, 43.30098, 40.51136, 40.51136, 40.51136, 
    40.51136, 40.51136, 40.51136, 40.51136, 40.51136, 40.51136, 40.51136, 
    40.51136, 40.51136, 40.51136, 40.51136, 40.51136, 40.51136, 40.51136, 
    40.51136, 40.51136, 40.51136, 40.51136, 40.51136, 40.51136, 40.51136, 
    40.51136, 40.51136, 40.51136, 40.51136, 40.51136, 40.51136, 40.51136, 
    40.51136, 40.51136, 40.51136, 40.51136, 40.51136, 40.51136, 40.22532,
  41.12221, 41.11818, 41.12221, 41.13429, 41.15435, 41.18228, 41.21794, 
    41.26115, 41.31168, 41.36928, 41.43365, 41.50449, 41.58142, 41.6641, 
    41.75211, 41.84505, 41.94248, 42.04395, 42.14902, 42.25722, 42.36808, 
    42.48113, 42.59591, 42.71193, 42.82874, 42.94588, 43.06289, 43.17934, 
    43.2948, 43.40885, 43.52108, 43.63111, 43.73857, 43.8431, 43.94437, 
    44.04205, 44.13586, 44.22551, 44.31076, 44.39137, 44.46712, 44.53784, 
    44.60335, 44.66352, 44.71823, 44.76739, 44.81092, 44.84879, 44.88097, 
    44.90746, 44.9283, 44.94352, 44.95322, 44.95747, 44.95641, 44.95018, 
    44.93893, 44.92284, 44.90213, 44.87702, 44.84774, 44.81456, 44.77774, 
    44.73758, 44.69438, 44.64846, 44.60015, 44.54979, 44.49771, 44.44429, 
    44.38987, 44.33482, 44.27951, 44.2243, 44.16957, 44.11565, 44.06293, 
    44.01173, 43.96241, 43.91528, 43.87065, 43.82883, 43.7901, 43.75471, 
    43.7229, 43.69488, 43.67084, 43.65095, 43.63534, 43.62411, 43.61734, 
    43.61508, 43.61734, 43.62411, 43.63534, 43.65095, 43.67084, 43.69488, 
    43.7229, 43.75471, 43.7901, 43.82883, 43.87065, 43.91528, 43.96241, 
    44.01173, 44.06293, 44.11565, 44.16957, 44.2243, 44.27951, 44.33482, 
    44.38987, 44.44429, 44.49771, 44.54979, 44.60015, 44.64846, 44.69438, 
    44.73758, 44.77774, 44.81456, 44.84774, 44.87702, 44.90213, 44.92284, 
    44.93893, 44.95018, 44.95641, 44.95747, 44.95322, 44.94352, 44.9283, 
    44.90746, 44.88097, 44.84879, 44.81092, 44.76739, 44.71823, 44.66352, 
    44.60335, 44.53784, 44.63784, 44.73784, 44.83784, 41.51136, 41.51136, 
    41.51136, 41.51136, 41.51136, 41.51136, 41.51136, 41.51136, 41.51136, 
    41.51136, 41.51136, 41.51136, 41.51136, 41.51136, 41.51136, 41.51136, 
    41.51136, 41.51136, 41.51136, 41.51136, 41.51136, 41.51136, 41.51136, 
    41.51136, 41.51136, 41.51136, 41.51136, 41.51136, 41.51136, 41.51136, 
    41.51136, 41.51136, 41.51136, 41.51136, 41.51136, 41.51136, 41.11818,
  41.94397, 41.93918, 41.94397, 41.95832, 41.98215, 42.01533, 42.05767, 
    42.10895, 42.1689, 42.23719, 42.31346, 42.39733, 42.48836, 42.5861, 
    42.69007, 42.79976, 42.91465, 43.03422, 43.1579, 43.28516, 43.41543, 
    43.54816, 43.68279, 43.81877, 43.95555, 44.09261, 44.22941, 44.36545, 
    44.50022, 44.63324, 44.76406, 44.89222, 45.01729, 45.13888, 45.2566, 
    45.37008, 45.479, 45.58302, 45.68187, 45.77529, 45.86303, 45.94487, 
    46.02064, 46.09018, 46.15335, 46.21006, 46.26022, 46.30378, 46.34073, 
    46.37107, 46.39483, 46.41208, 46.42289, 46.42738, 46.4257, 46.418, 
    46.40447, 46.38533, 46.3608, 46.33115, 46.29666, 46.25762, 46.21435, 
    46.16718, 46.11647, 46.06258, 46.00589, 45.9468, 45.88571, 45.82303, 
    45.75918, 45.69458, 45.62966, 45.56484, 45.50056, 45.43724, 45.37528, 
    45.31511, 45.25712, 45.20169, 45.1492, 45.09999, 45.0544, 45.01273, 
    44.97527, 44.94226, 44.91394, 44.8905, 44.8721, 44.85886, 44.85089, 
    44.84822, 44.85089, 44.85886, 44.8721, 44.8905, 44.91394, 44.94226, 
    44.97527, 45.01273, 45.0544, 45.09999, 45.1492, 45.20169, 45.25712, 
    45.31511, 45.37528, 45.43724, 45.50056, 45.56484, 45.62966, 45.69458, 
    45.75918, 45.82303, 45.88571, 45.9468, 46.00589, 46.06258, 46.11647, 
    46.16718, 46.21435, 46.25762, 46.29666, 46.33115, 46.3608, 46.38533, 
    46.40447, 46.418, 46.4257, 46.42738, 46.42289, 46.41208, 46.39483, 
    46.37107, 46.34073, 46.30378, 46.26022, 46.21006, 46.15335, 46.09018, 
    46.02064, 45.94487, 46.04487, 46.14487, 46.24487, 46.34487, 42.51136, 
    42.51136, 42.51136, 42.51136, 42.51136, 42.51136, 42.51136, 42.51136, 
    42.51136, 42.51136, 42.51136, 42.51136, 42.51136, 42.51136, 42.51136, 
    42.51136, 42.51136, 42.51136, 42.51136, 42.51136, 42.51136, 42.51136, 
    42.51136, 42.51136, 42.51136, 42.51136, 42.51136, 42.51136, 42.51136, 
    42.51136, 42.51136, 42.51136, 42.51136, 42.51136, 42.51136, 41.93918,
  42.69794, 42.69231, 42.69794, 42.71479, 42.74277, 42.78172, 42.83141, 
    42.89155, 42.96182, 43.04181, 43.1311, 43.22919, 43.33558, 43.4497, 
    43.57098, 43.69882, 43.83259, 43.97166, 44.11539, 44.26311, 44.41419, 
    44.56797, 44.72381, 44.88106, 45.0391, 45.19731, 45.35509, 45.51186, 
    45.66705, 45.82011, 45.97052, 46.11776, 46.26137, 46.40088, 46.53585, 
    46.6659, 46.79062, 46.90968, 47.02275, 47.12952, 47.22975, 47.32318, 
    47.40961, 47.48887, 47.56081, 47.62532, 47.6823, 47.73172, 47.77354, 
    47.80778, 47.83447, 47.85369, 47.86553, 47.87012, 47.86764, 47.85825, 
    47.84218, 47.81967, 47.79099, 47.75642, 47.71629, 47.67094, 47.62073, 
    47.56604, 47.50727, 47.44484, 47.37919, 47.31076, 47.24002, 47.16744, 
    47.09349, 47.01867, 46.94347, 46.86837, 46.79387, 46.72045, 46.64861, 
    46.57881, 46.51152, 46.44719, 46.38624, 46.32908, 46.27612, 46.22769, 
    46.18414, 46.14576, 46.11282, 46.08556, 46.06415, 46.04875, 46.03947, 
    46.03637, 46.03947, 46.04875, 46.06415, 46.08556, 46.11282, 46.14576, 
    46.18414, 46.22769, 46.27612, 46.32908, 46.38624, 46.44719, 46.51152, 
    46.57881, 46.64861, 46.72045, 46.79387, 46.86837, 46.94347, 47.01867, 
    47.09349, 47.16744, 47.24002, 47.31076, 47.37919, 47.44484, 47.50727, 
    47.56604, 47.62073, 47.67094, 47.71629, 47.75642, 47.79099, 47.81967, 
    47.84218, 47.85825, 47.86764, 47.87012, 47.86553, 47.85369, 47.83447, 
    47.80778, 47.77354, 47.73172, 47.6823, 47.62532, 47.56081, 47.48887, 
    47.40961, 47.32318, 47.42318, 47.52318, 47.62318, 47.72318, 43.51136, 
    43.51136, 43.51136, 43.51136, 43.51136, 43.51136, 43.51136, 43.51136, 
    43.51136, 43.51136, 43.51136, 43.51136, 43.51136, 43.51136, 43.51136, 
    43.51136, 43.51136, 43.51136, 43.51136, 43.51136, 43.51136, 43.51136, 
    43.51136, 43.51136, 43.51136, 43.51136, 43.51136, 43.51136, 43.51136, 
    43.51136, 43.51136, 43.51136, 43.51136, 43.51136, 43.51136, 42.69231,
  43.38826, 43.38171, 43.38826, 43.40785, 43.44038, 43.48565, 43.54336, 
    43.61319, 43.6947, 43.78744, 43.89085, 44.00437, 44.12737, 44.25918, 
    44.39911, 44.54644, 44.70045, 44.86039, 45.02549, 45.19501, 45.3682, 
    45.5443, 45.72256, 45.90227, 46.08271, 46.26317, 46.44299, 46.6215, 
    46.79806, 46.97207, 47.14293, 47.31008, 47.47298, 47.63114, 47.78405, 
    47.93128, 48.07241, 48.20704, 48.33481, 48.4554, 48.56852, 48.67389, 
    48.77131, 48.86056, 48.94149, 49.01397, 49.07792, 49.13328, 49.18002, 
    49.21816, 49.24775, 49.26886, 49.2816, 49.28614, 49.28265, 49.27134, 
    49.25245, 49.22625, 49.19306, 49.1532, 49.10703, 49.05492, 48.9973, 
    48.9346, 48.86726, 48.79575, 48.72058, 48.64223, 48.56125, 48.47816, 
    48.3935, 48.30783, 48.22171, 48.13569, 48.05033, 47.96621, 47.88385, 
    47.80381, 47.72663, 47.65281, 47.58285, 47.51723, 47.45639, 47.40075, 
    47.3507, 47.30658, 47.26871, 47.23735, 47.21273, 47.19501, 47.18433, 
    47.18077, 47.18433, 47.19501, 47.21273, 47.23735, 47.26871, 47.30658, 
    47.3507, 47.40075, 47.45639, 47.51723, 47.58285, 47.65281, 47.72663, 
    47.80381, 47.88385, 47.96621, 48.05033, 48.13569, 48.22171, 48.30783, 
    48.3935, 48.47816, 48.56125, 48.64223, 48.72058, 48.79575, 48.86726, 
    48.9346, 48.9973, 49.05492, 49.10703, 49.1532, 49.19306, 49.22625, 
    49.25245, 49.27134, 49.28265, 49.28614, 49.2816, 49.26886, 49.24775, 
    49.21816, 49.18002, 49.13328, 49.07792, 49.01397, 48.94149, 48.86056, 
    48.77131, 48.67389, 48.7739, 48.87389, 48.97389, 49.07389, 44.51136, 
    44.51136, 44.51136, 44.51136, 44.51136, 44.51136, 44.51136, 44.51136, 
    44.51136, 44.51136, 44.51136, 44.51136, 44.51136, 44.51136, 44.51136, 
    44.51136, 44.51136, 44.51136, 44.51136, 44.51136, 44.51136, 44.51136, 
    44.51136, 44.51136, 44.51136, 44.51136, 44.51136, 44.51136, 44.51136, 
    44.51136, 44.51136, 44.51136, 44.51136, 44.51136, 44.51136, 43.38171,
  44.01912, 44.01157, 44.01912, 44.04171, 44.0792, 44.13135, 44.19781, 
    44.27816, 44.37188, 44.47841, 44.5971, 44.72725, 44.86811, 45.01889, 
    45.17877, 45.34691, 45.52246, 45.70454, 45.89228, 46.08482, 46.2813, 
    46.48085, 46.68264, 46.88586, 47.08969, 47.29337, 47.49612, 47.69723, 
    47.89598, 48.09169, 48.28373, 48.47146, 48.65429, 48.83168, 49.00308, 
    49.16801, 49.326, 49.47663, 49.6195, 49.75426, 49.88057, 49.99817, 
    50.10679, 50.20623, 50.29631, 50.37689, 50.44788, 50.50922, 50.56088, 
    50.60288, 50.63528, 50.65816, 50.67167, 50.67596, 50.67123, 50.65773, 
    50.63573, 50.60554, 50.56749, 50.52195, 50.46933, 50.41005, 50.34457, 
    50.27337, 50.19696, 50.11586, 50.03063, 49.94183, 49.85005, 49.75588, 
    49.65994, 49.56284, 49.46521, 49.36768, 49.27088, 49.17545, 49.082, 
    48.99116, 48.90352, 48.81968, 48.74019, 48.66561, 48.59644, 48.53316, 
    48.47622, 48.42602, 48.38291, 48.34721, 48.31917, 48.29899, 48.28683, 
    48.28276, 48.28683, 48.29899, 48.31917, 48.34721, 48.38291, 48.42602, 
    48.47622, 48.53316, 48.59644, 48.66561, 48.74019, 48.81968, 48.90352, 
    48.99116, 49.082, 49.17545, 49.27088, 49.36768, 49.46521, 49.56284, 
    49.65994, 49.75588, 49.85005, 49.94183, 50.03063, 50.11586, 50.19696, 
    50.27337, 50.34457, 50.41005, 50.46933, 50.52195, 50.56749, 50.60554, 
    50.63573, 50.65773, 50.67123, 50.67596, 50.67167, 50.65816, 50.63528, 
    50.60288, 50.56088, 50.50922, 50.44788, 50.37689, 50.29631, 50.20623, 
    50.10679, 49.99817, 50.09817, 50.19817, 50.29817, 50.39817, 45.51136, 
    45.51136, 45.51136, 45.51136, 45.51136, 45.51136, 45.51136, 45.51136, 
    45.51136, 45.51136, 45.51136, 45.51136, 45.51136, 45.51136, 45.51136, 
    45.51136, 45.51136, 45.51136, 45.51136, 45.51136, 45.51136, 45.51136, 
    45.51136, 45.51136, 45.51136, 45.51136, 45.51136, 45.51136, 45.51136, 
    45.51136, 45.51136, 45.51136, 45.51136, 45.51136, 45.51136, 44.01157,
  44.5947, 44.58606, 44.5947, 44.62056, 44.66346, 44.72308, 44.79903, 
    44.89077, 44.9977, 45.11911, 45.25423, 45.40221, 45.56218, 45.73318, 
    45.91428, 46.10448, 46.3028, 46.50822, 46.71976, 46.93643, 47.15726, 
    47.38128, 47.60757, 47.83519, 48.06328, 48.29097, 48.51741, 48.74182, 
    48.96342, 49.18146, 49.39524, 49.60409, 49.80735, 50.00443, 50.19475, 
    50.37777, 50.55299, 50.71995, 50.87822, 51.0274, 51.16715, 51.29716, 
    51.41716, 51.52691, 51.62624, 51.71497, 51.79303, 51.86034, 51.91687, 
    51.96265, 51.99775, 52.02227, 52.03634, 52.04017, 52.03397, 52.01801, 
    51.9926, 51.95807, 51.9148, 51.86321, 51.80373, 51.73685, 51.66307, 
    51.58292, 51.49696, 51.40578, 51.31, 51.21023, 51.10712, 51.00135, 
    50.89358, 50.78451, 50.67483, 50.56525, 50.45646, 50.34919, 50.24411, 
    50.14193, 50.04333, 49.94896, 49.85947, 49.77546, 49.69753, 49.62621, 
    49.56201, 49.50539, 49.45676, 49.41648, 49.38484, 49.36206, 49.34833, 
    49.34374, 49.34833, 49.36206, 49.38484, 49.41648, 49.45676, 49.50539, 
    49.56201, 49.62621, 49.69753, 49.77546, 49.85947, 49.94896, 50.04333, 
    50.14193, 50.24411, 50.34919, 50.45646, 50.56525, 50.67483, 50.78451, 
    50.89358, 51.00135, 51.10712, 51.21023, 51.31, 51.40578, 51.49696, 
    51.58292, 51.66307, 51.73685, 51.80373, 51.86321, 51.9148, 51.95807, 
    51.9926, 52.01801, 52.03397, 52.04017, 52.03634, 52.02227, 51.99775, 
    51.96265, 51.91687, 51.86034, 51.79303, 51.71497, 51.62624, 51.52691, 
    51.41716, 51.29716, 51.16715, 51.0274, 50.87822, 50.71995, 50.55299, 
    50.37777, 50.19475, 50.00443, 49.80735, 49.60409, 49.39524, 49.18146, 
    48.96342, 48.74182, 48.51741, 48.29097, 48.06328, 47.83519, 47.60757, 
    47.38128, 46.51136, 46.51136, 46.51136, 46.51136, 46.51136, 46.51136, 
    46.51136, 46.51136, 46.51136, 46.51136, 46.51136, 46.51136, 46.51136, 
    46.51136, 46.51136, 46.51136, 46.51136, 46.51136, 46.51136, 44.58606,
  45.11909, 45.10926, 45.11909, 45.14849, 45.19726, 45.265, 45.35122, 
    45.45528, 45.57643, 45.71383, 45.86655, 46.03358, 46.21389, 46.40636, 
    46.6099, 46.82335, 47.04558, 47.27545, 47.51184, 47.75363, 47.99974, 
    48.24911, 48.50069, 48.75349, 49.00654, 49.25888, 49.50962, 49.75789, 
    50.00285, 50.2437, 50.47967, 50.71004, 50.93412, 51.15124, 51.36079, 
    51.5622, 51.75492, 51.93844, 52.11232, 52.27612, 52.42946, 52.57202, 
    52.70349, 52.82363, 52.93224, 53.02915, 53.11425, 53.18747, 53.2488, 
    53.29825, 53.3359, 53.36187, 53.37631, 53.37944, 53.3715, 53.35279, 
    53.32364, 53.28444, 53.2356, 53.17756, 53.11083, 53.03592, 52.9534, 
    52.86385, 52.76789, 52.66617, 52.55935, 52.44812, 52.3332, 52.21532, 
    52.09523, 51.97369, 51.85145, 51.72931, 51.60804, 51.48842, 51.37123, 
    51.25723, 51.14719, 51.04184, 50.94189, 50.84804, 50.76094, 50.6812, 
    50.60941, 50.54607, 50.49165, 50.44656, 50.41114, 50.38564, 50.37026, 
    50.36512, 50.37026, 50.38564, 50.41114, 50.44656, 50.49165, 50.54607, 
    50.60941, 50.6812, 50.76094, 50.84804, 50.94189, 51.04184, 51.14719, 
    51.25723, 51.37123, 51.48842, 51.60804, 51.72931, 51.85145, 51.97369, 
    52.09523, 52.21532, 52.3332, 52.44812, 52.55935, 52.66617, 52.76789, 
    52.86385, 52.9534, 53.03592, 53.11083, 53.17756, 53.2356, 53.28444, 
    53.32364, 53.35279, 53.3715, 53.37944, 53.37631, 53.36187, 53.3359, 
    53.29825, 53.2488, 53.18747, 53.11425, 53.02915, 52.93224, 52.82363, 
    52.70349, 52.57202, 52.42946, 52.27612, 52.11232, 51.93844, 51.75492, 
    51.5622, 51.36079, 51.15124, 50.93412, 50.71004, 50.47967, 50.2437, 
    50.00285, 49.75789, 49.50962, 49.25888, 49.00654, 48.75349, 48.50069, 
    48.24911, 47.51136, 47.51136, 47.51136, 47.51136, 47.51136, 47.51136, 
    47.51136, 47.51136, 47.51136, 47.51136, 47.51136, 47.51136, 47.51136, 
    47.51136, 47.51136, 47.51136, 47.51136, 47.51136, 47.51136, 45.10926,
  45.59623, 45.58511, 45.59623, 45.62949, 45.68462, 45.76115, 45.85847, 
    45.97581, 46.11226, 46.26679, 46.4383, 46.62561, 46.82747, 47.04261, 
    47.26974, 47.50756, 47.75477, 48.01009, 48.27225, 48.54003, 48.81222, 
    49.08765, 49.3652, 49.64378, 49.92233, 50.19983, 50.47532, 50.74787, 
    51.01657, 51.28057, 51.53905, 51.79123, 52.03638, 52.2738, 52.50281, 
    52.72281, 52.9332, 53.13346, 53.32309, 53.50163, 53.66867, 53.82385, 
    53.96685, 54.09742, 54.21531, 54.32037, 54.41246, 54.49152, 54.55753, 
    54.61051, 54.65054, 54.67775, 54.69233, 54.6945, 54.68454, 54.66277, 
    54.62955, 54.58532, 54.53052, 54.46566, 54.39126, 54.30791, 54.21622, 
    54.11683, 54.01041, 53.89769, 53.77937, 53.65622, 53.52903, 53.39858, 
    53.2657, 53.13121, 52.99597, 52.86081, 52.72659, 52.59417, 52.46442, 
    52.33816, 52.21624, 52.09948, 51.98868, 51.88459, 51.78796, 51.69946, 
    51.61975, 51.54941, 51.48896, 51.43885, 51.39948, 51.37114, 51.35404, 
    51.34833, 51.35404, 51.37114, 51.39948, 51.43885, 51.48896, 51.54941, 
    51.61975, 51.69946, 51.78796, 51.88459, 51.98868, 52.09948, 52.21624, 
    52.33816, 52.46442, 52.59417, 52.72659, 52.86081, 52.99597, 53.13121, 
    53.2657, 53.39858, 53.52903, 53.65622, 53.77937, 53.89769, 54.01041, 
    54.11683, 54.21622, 54.30791, 54.39126, 54.46566, 54.53052, 54.58532, 
    54.62955, 54.66277, 54.68454, 54.6945, 54.69233, 54.67775, 54.65054, 
    54.61051, 54.55753, 54.49152, 54.41246, 54.32037, 54.21531, 54.09742, 
    53.96685, 53.82385, 53.66867, 53.50163, 53.32309, 53.13346, 52.9332, 
    52.72281, 52.50281, 52.2738, 52.03638, 51.79123, 51.53905, 51.28057, 
    51.01657, 50.74787, 50.47532, 50.19983, 49.92233, 49.64378, 49.3652, 
    49.08765, 48.81222, 48.54003, 48.27225, 48.01009, 47.75477, 47.50756, 
    47.26974, 47.04261, 46.82747, 46.62561, 46.4383, 46.26679, 46.11226, 
    45.97581, 45.85847, 45.76115, 45.68462, 45.62949, 45.59623, 45.58511,
  46.02989, 46.01737, 46.02989, 46.06734, 46.12937, 46.21543, 46.32474, 
    46.45637, 46.60922, 46.78206, 46.97358, 47.18237, 47.40699, 47.64595, 
    47.89779, 48.161, 48.43415, 48.71579, 49.00453, 49.29901, 49.59792, 49.9, 
    50.20403, 50.50883, 50.81328, 51.1163, 51.41686, 51.71395, 52.00665, 
    52.29402, 52.57521, 52.8494, 53.1158, 53.37366, 53.62228, 53.861, 
    54.08919, 54.30629, 54.51176, 54.70511, 54.88591, 55.05375, 55.20831, 
    55.34929, 55.47644, 55.58959, 55.6886, 55.77339, 55.84394, 55.90028, 
    55.9425, 55.97074, 55.9852, 55.98614, 55.97384, 55.94868, 55.91106, 
    55.86142, 55.80029, 55.72818, 55.64571, 55.55349, 55.45219, 55.34253, 
    55.22522, 55.10104, 54.97078, 54.83527, 54.69535, 54.5519, 54.4058, 
    54.25794, 54.10925, 53.96064, 53.81306, 53.66744, 53.52471, 53.3858, 
    53.25162, 53.12308, 53.00104, 52.88637, 52.77987, 52.6823, 52.59438, 
    52.51677, 52.45006, 52.39474, 52.35126, 52.31996, 52.30108, 52.29477, 
    52.30108, 52.31996, 52.35126, 52.39474, 52.45006, 52.51677, 52.59438, 
    52.6823, 52.77987, 52.88637, 53.00104, 53.12308, 53.25162, 53.3858, 
    53.52471, 53.66744, 53.81306, 53.96064, 54.10925, 54.25794, 54.4058, 
    54.5519, 54.69535, 54.83527, 54.97078, 55.10104, 55.22522, 55.34253, 
    55.45219, 55.55349, 55.64571, 55.72818, 55.80029, 55.86142, 55.91106, 
    55.94868, 55.97384, 55.98614, 55.9852, 55.97074, 55.9425, 55.90028, 
    55.84394, 55.77339, 55.6886, 55.58959, 55.47644, 55.34929, 55.20831, 
    55.05375, 54.88591, 54.70511, 54.51176, 54.30629, 54.08919, 53.861, 
    53.62228, 53.37366, 53.1158, 52.8494, 52.57521, 52.29402, 52.00665, 
    51.71395, 51.41686, 51.1163, 50.81328, 50.50883, 50.20403, 49.9, 
    49.59792, 49.29901, 49.00453, 48.71579, 48.43415, 48.161, 47.89779, 
    47.64595, 47.40699, 47.18237, 46.97358, 46.78206, 46.60922, 46.45637, 
    46.32474, 46.21543, 46.12937, 46.06734, 46.02989, 46.01737,
  46.42366, 46.40962, 46.42366, 46.46566, 46.53519, 46.63155, 46.7538, 
    46.9008, 47.07122, 47.26359, 47.47634, 47.70782, 47.95636, 48.22025, 
    48.4978, 48.78735, 49.08727, 49.39598, 49.71195, 50.03371, 50.35984, 
    50.68898, 51.01984, 51.35117, 51.68178, 52.01052, 52.33632, 52.65813, 
    52.97495, 53.28581, 53.58982, 53.88611, 54.17384, 54.45223, 54.72053, 
    54.97804, 55.2241, 55.4581, 55.67947, 55.88767, 56.08225, 56.26278, 
    56.42889, 56.58026, 56.71663, 56.83781, 56.94363, 57.03403, 57.10897, 
    57.16849, 57.21268, 57.24171, 57.25578, 57.25518, 57.24024, 57.21134, 
    57.16893, 57.11351, 57.04562, 56.96587, 56.87489, 56.77337, 56.66203, 
    56.54164, 56.41299, 56.27692, 56.13429, 55.98599, 55.83293, 55.67605, 
    55.51631, 55.35468, 55.19215, 55.02972, 54.8684, 54.7092, 54.55313, 
    54.40121, 54.25442, 54.11375, 53.98016, 53.85458, 53.73791, 53.63099, 
    53.5346, 53.44949, 53.3763, 53.3156, 53.26788, 53.23351, 53.21278, 
    53.20585, 53.21278, 53.23351, 53.26788, 53.3156, 53.3763, 53.44949, 
    53.5346, 53.63099, 53.73791, 53.85458, 53.98016, 54.11375, 54.25442, 
    54.40121, 54.55313, 54.7092, 54.8684, 55.02972, 55.19215, 55.35468, 
    55.51631, 55.67605, 55.83293, 55.98599, 56.13429, 56.27692, 56.41299, 
    56.54164, 56.66203, 56.77337, 56.87489, 56.96587, 57.04562, 57.11351, 
    57.16893, 57.21134, 57.24024, 57.25518, 57.25578, 57.24171, 57.21268, 
    57.16849, 57.10897, 57.03403, 56.94363, 56.83781, 56.71663, 56.58026, 
    56.42889, 56.26278, 56.08225, 55.88767, 55.67947, 55.4581, 55.2241, 
    54.97804, 54.72053, 54.45223, 54.17384, 53.88611, 53.58982, 53.28581, 
    52.97495, 52.65813, 52.33632, 52.01052, 51.68178, 51.35117, 51.01984, 
    50.68898, 50.35984, 50.03371, 49.71195, 49.39598, 49.08727, 48.78735, 
    48.4978, 48.22025, 47.95636, 47.70782, 47.47634, 47.26359, 47.07122, 
    46.9008, 46.7538, 46.63155, 46.53519, 46.46566, 46.42366, 46.40962,
  46.78093, 46.76522, 46.78093, 46.82788, 46.90554, 47.01306, 47.14927, 
    47.31279, 47.50199, 47.71513, 47.95034, 48.20571, 48.47929, 48.76913, 
    49.07333, 49.39003, 49.71744, 50.05383, 50.39754, 50.74698, 51.10066, 
    51.45713, 51.81502, 52.17303, 52.52991, 52.88446, 53.23556, 53.58212, 
    53.92308, 54.25747, 54.58431, 54.90271, 55.2118, 55.51074, 55.79875, 
    56.07509, 56.33905, 56.58998, 56.82727, 57.05036, 57.25874, 57.45195, 
    57.62959, 57.79132, 57.93686, 58.06598, 58.17852, 58.27439, 58.35356, 
    58.41607, 58.46201, 58.49156, 58.50496, 58.50251, 58.48457, 58.45156, 
    58.40398, 58.34237, 58.26731, 58.17947, 58.07954, 57.96827, 57.84643, 
    57.71487, 57.57444, 57.42604, 57.2706, 57.10909, 56.94247, 56.77177, 
    56.59801, 56.42224, 56.24551, 56.0689, 55.8935, 55.72039, 55.55066, 
    55.38541, 55.2257, 55.07261, 54.92718, 54.79042, 54.66331, 54.54678, 
    54.44169, 54.34886, 54.269, 54.20276, 54.15067, 54.11314, 54.0905, 
    54.08293, 54.0905, 54.11314, 54.15067, 54.20276, 54.269, 54.34886, 
    54.44169, 54.54678, 54.66331, 54.79042, 54.92718, 55.07261, 55.2257, 
    55.38541, 55.55066, 55.72039, 55.8935, 56.0689, 56.24551, 56.42224, 
    56.59801, 56.77177, 56.94247, 57.10909, 57.2706, 57.42604, 57.57444, 
    57.71487, 57.84643, 57.96827, 58.07954, 58.17947, 58.26731, 58.34237, 
    58.40398, 58.45156, 58.48457, 58.50251, 58.50496, 58.49156, 58.46201, 
    58.41607, 58.35356, 58.27439, 58.17852, 58.06598, 57.93686, 57.79132, 
    57.62959, 57.45195, 57.25874, 57.05036, 56.82727, 56.58998, 56.33905, 
    56.07509, 55.79875, 55.51074, 55.2118, 54.90271, 54.58431, 54.25747, 
    53.92308, 53.58212, 53.23556, 52.88446, 52.52991, 52.17303, 51.81502, 
    51.45713, 51.10066, 50.74698, 50.39754, 50.05383, 49.71744, 49.39003, 
    49.07333, 48.76913, 48.47929, 48.20571, 47.95034, 47.71513, 47.50199, 
    47.31279, 47.14927, 47.01306, 46.90554, 46.82788, 46.78093, 46.76522,
  47.10486, 47.08733, 47.10486, 47.1572, 47.24371, 47.36332, 47.5146, 
    47.69584, 47.9051, 48.14029, 48.3992, 48.67961, 48.97927, 49.29601, 
    49.62767, 49.97221, 50.32767, 50.69219, 51.06398, 51.44137, 51.82277, 
    52.20667, 52.59165, 52.97635, 53.35948, 53.7398, 54.11614, 54.48738, 
    54.85244, 55.21027, 55.55991, 55.90038, 56.2308, 56.55027, 56.85799, 
    57.15316, 57.43503, 57.70291, 57.95614, 58.19413, 58.41632, 58.62222, 
    58.81139, 58.98345, 59.1381, 59.27509, 59.39425, 59.49545, 59.57868, 
    59.64397, 59.69143, 59.72124, 59.73366, 59.72902, 59.70772, 59.67022, 
    59.61705, 59.54881, 59.46614, 59.36975, 59.26041, 59.13891, 59.00611, 
    58.86292, 58.71025, 58.54908, 58.38041, 58.20526, 58.02469, 57.83978, 
    57.65163, 57.46136, 57.2701, 57.07899, 56.88921, 56.70189, 56.51823, 
    56.33937, 56.16648, 56.00071, 55.84319, 55.69501, 55.55723, 55.43087, 
    55.31688, 55.21615, 55.12946, 55.05753, 55.00095, 54.96018, 54.93558, 
    54.92736, 54.93558, 54.96018, 55.00095, 55.05753, 55.12946, 55.21615, 
    55.31688, 55.43087, 55.55723, 55.69501, 55.84319, 56.00071, 56.16648, 
    56.33937, 56.51823, 56.70189, 56.88921, 57.07899, 57.2701, 57.46136, 
    57.65163, 57.83978, 58.02469, 58.20526, 58.38041, 58.54908, 58.71025, 
    58.86292, 59.00611, 59.13891, 59.26041, 59.36975, 59.46614, 59.54881, 
    59.61705, 59.67022, 59.70772, 59.72902, 59.73366, 59.72124, 59.69143, 
    59.64397, 59.57868, 59.49545, 59.39425, 59.27509, 59.1381, 58.98345, 
    58.81139, 58.62222, 58.41632, 58.19413, 57.95614, 57.70291, 57.43503, 
    57.15316, 56.85799, 56.55027, 56.2308, 55.90038, 55.55991, 55.21027, 
    54.85244, 54.48738, 54.11614, 53.7398, 53.35948, 52.97635, 52.59165, 
    52.20667, 51.82277, 51.44137, 51.06398, 50.69219, 50.32767, 49.97221, 
    49.62767, 49.29601, 48.97927, 48.67961, 48.3992, 48.14029, 47.9051, 
    47.69584, 47.5146, 47.36332, 47.24371, 47.1572, 47.10486, 47.08733,
  47.3984, 47.37889, 47.3984, 47.45664, 47.55278, 47.6855, 47.85304, 48.0533, 
    48.28394, 48.54247, 48.82631, 49.13286, 49.45959, 49.80405, 50.16385, 
    50.53677, 50.92068, 51.31361, 51.71366, 52.11908, 52.52822, 52.93951, 
    53.35149, 53.76276, 54.172, 54.57793, 54.97937, 55.37514, 55.76414, 
    56.14531, 56.51762, 56.88009, 57.23177, 57.57174, 57.89913, 58.21312, 
    58.51291, 58.79776, 59.06696, 59.31987, 59.5559, 59.7745, 59.9752, 
    60.15759, 60.32131, 60.46611, 60.59177, 60.69819, 60.78531, 60.85318, 
    60.90191, 60.9317, 60.94283, 60.93565, 60.9106, 60.86819, 60.80899, 
    60.73366, 60.6429, 60.53748, 60.41823, 60.28602, 60.14177, 59.98646, 
    59.82109, 59.64669, 59.46434, 59.27515, 59.08023, 58.88074, 58.67786, 
    58.47276, 58.26665, 58.06076, 57.85631, 57.65454, 57.45669, 57.264, 
    57.07772, 56.89906, 56.72924, 56.56944, 56.4208, 56.28443, 56.16137, 
    56.05257, 55.95891, 55.88117, 55.82, 55.77592, 55.74932, 55.74042, 
    55.74932, 55.77592, 55.82, 55.88117, 55.95891, 56.05257, 56.16137, 
    56.28443, 56.4208, 56.56944, 56.72924, 56.89906, 57.07772, 57.264, 
    57.45669, 57.65454, 57.85631, 58.06076, 58.26665, 58.47276, 58.67786, 
    58.88074, 59.08023, 59.27515, 59.46434, 59.64669, 59.82109, 59.98646, 
    60.14177, 60.28602, 60.41823, 60.53748, 60.6429, 60.73366, 60.80899, 
    60.86819, 60.9106, 60.93565, 60.94283, 60.9317, 60.90191, 60.85318, 
    60.78531, 60.69819, 60.59177, 60.46611, 60.32131, 60.15759, 59.9752, 
    59.7745, 59.5559, 59.31987, 59.06696, 58.79776, 58.51291, 58.21312, 
    57.89913, 57.57174, 57.23177, 56.88009, 56.51762, 56.14531, 55.76414, 
    55.37514, 54.97937, 54.57793, 54.172, 53.76276, 53.35149, 52.93951, 
    52.52822, 52.11908, 51.71366, 51.31361, 50.92068, 50.53677, 50.16385, 
    49.80405, 49.45959, 49.13286, 48.82631, 48.54247, 48.28394, 48.0533, 
    47.85304, 47.6855, 47.55278, 47.45664, 47.3984, 47.37889,
  47.6643, 47.64262, 47.6643, 47.72899, 47.83565, 47.98261, 48.1677, 
    48.38836, 48.64175, 48.92492, 49.23486, 49.56859, 49.92326, 50.29612, 
    50.68459, 51.08626, 51.49886, 51.9203, 52.34861, 52.78199, 53.21873, 
    53.65722, 54.09598, 54.53358, 54.96867, 55.39997, 55.82625, 56.24634, 
    56.65909, 57.06342, 57.45827, 57.84261, 58.21546, 58.57586, 58.92291, 
    59.25571, 59.57344, 59.87529, 60.1605, 60.42839, 60.6783, 60.90965, 
    61.1219, 61.31462, 61.4874, 61.63996, 61.77206, 61.88357, 61.97443, 
    62.04467, 62.09443, 62.12391, 62.1334, 62.12331, 62.09411, 62.04635, 
    61.98066, 61.89775, 61.79839, 61.68341, 61.55373, 61.41028, 61.25407, 
    61.08614, 60.90757, 60.71947, 60.52301, 60.31935, 60.10969, 59.89526, 
    59.6773, 59.45706, 59.23583, 59.01489, 58.79555, 58.5791, 58.36686, 
    58.16016, 57.96029, 57.76857, 57.5863, 57.41472, 57.25508, 57.10855, 
    56.97628, 56.85929, 56.75854, 56.67489, 56.60905, 56.5616, 56.53295, 
    56.52337, 56.53295, 56.5616, 56.60905, 56.67489, 56.75854, 56.85929, 
    56.97628, 57.10855, 57.25508, 57.41472, 57.5863, 57.76857, 57.96029, 
    58.16016, 58.36686, 58.5791, 58.79555, 59.01489, 59.23583, 59.45706, 
    59.6773, 59.89526, 60.10969, 60.31935, 60.52301, 60.71947, 60.90757, 
    61.08614, 61.25407, 61.41028, 61.55373, 61.68341, 61.79839, 61.89775, 
    61.98066, 62.04635, 62.09411, 62.12331, 62.1334, 62.12391, 62.09443, 
    62.04467, 61.97443, 61.88357, 61.77206, 61.63996, 61.4874, 61.31462, 
    61.1219, 60.90965, 60.6783, 60.42839, 60.1605, 59.87529, 59.57344, 
    59.25571, 58.92291, 58.57586, 58.21546, 57.84261, 57.45827, 57.06342, 
    56.65909, 56.24634, 55.82625, 55.39997, 54.96867, 54.53358, 54.09598, 
    53.65722, 53.21873, 52.78199, 52.34861, 51.9203, 51.49886, 51.08626, 
    50.68459, 50.29612, 49.92326, 49.56859, 49.23486, 48.92492, 48.64175, 
    48.38836, 48.1677, 47.98261, 47.83565, 47.72899, 47.6643, 47.64262,
  47.90511, 47.88103, 47.90511, 47.97689, 48.09505, 48.2575, 48.46154, 
    48.70403, 48.98157, 49.29067, 49.62783, 49.98968, 50.37301, 50.77482, 
    51.19231, 51.6229, 52.06423, 52.51411, 52.97053, 53.43163, 53.89566, 
    54.36104, 54.82623, 55.28979, 55.7504, 56.20673, 56.65755, 57.10167, 
    57.53793, 57.96521, 58.38241, 58.7885, 59.18243, 59.56322, 59.9299, 
    60.28153, 60.61723, 60.93614, 61.23744, 61.52039, 61.78427, 62.02844, 
    62.25232, 62.45541, 62.63728, 62.79758, 62.93607, 63.05256, 63.14701, 
    63.21943, 63.26996, 63.29883, 63.30635, 63.29296, 63.25916, 63.20558, 
    63.13288, 63.04187, 62.93336, 62.80828, 62.6676, 62.51236, 62.34363, 
    62.16255, 61.97027, 61.76799, 61.55695, 61.33839, 61.1136, 60.88386, 
    60.65049, 60.41483, 60.17822, 59.942, 59.70755, 59.47624, 59.24946, 
    59.02859, 58.81502, 58.61012, 58.41527, 58.23181, 58.06106, 57.90428, 
    57.76269, 57.63742, 57.5295, 57.43986, 57.36929, 57.31841, 57.28769, 
    57.27742, 57.28769, 57.31841, 57.36929, 57.43986, 57.5295, 57.63742, 
    57.76269, 57.90428, 58.06106, 58.23181, 58.41527, 58.61012, 58.81502, 
    59.02859, 59.24946, 59.47624, 59.70755, 59.942, 60.17822, 60.41483, 
    60.65049, 60.88386, 61.1136, 61.33839, 61.55695, 61.76799, 61.97027, 
    62.16255, 62.34363, 62.51236, 62.6676, 62.80828, 62.93336, 63.04187, 
    63.13288, 63.20558, 63.25916, 63.29296, 63.30635, 63.29883, 63.26996, 
    63.21943, 63.14701, 63.05256, 62.93607, 62.79758, 62.63728, 62.45541, 
    62.25232, 62.02844, 61.78427, 61.52039, 61.23744, 60.93614, 60.61723, 
    60.28153, 59.9299, 59.56322, 59.18243, 58.7885, 58.38241, 57.96521, 
    57.53793, 57.10167, 56.65755, 56.20673, 55.7504, 55.28979, 54.82623, 
    54.36104, 53.89566, 53.43163, 52.97053, 52.51411, 52.06423, 51.6229, 
    51.19231, 50.77482, 50.37301, 49.98968, 49.62783, 49.29067, 48.98157, 
    48.70403, 48.46154, 48.2575, 48.09505, 47.97689, 47.90511, 47.88103,
  48.12318, 48.09645, 48.12318, 48.20277, 48.33353, 48.51285, 48.73734, 
    49.00319, 49.3063, 49.64257, 50.00798, 50.39874, 50.8113, 51.2424, 
    51.68906, 52.14857, 52.61848, 53.09655, 53.58073, 54.06915, 54.56006, 
    55.05185, 55.54301, 56.03211, 56.51779, 56.99876, 57.47375, 57.94158, 
    58.40106, 58.85105, 59.29044, 59.71813, 60.13306, 60.53419, 60.9205, 
    61.291, 61.64475, 61.98082, 62.29833, 62.59647, 62.87445, 63.13157, 
    63.3672, 63.58075, 63.77176, 63.93984, 64.08468, 64.20609, 64.304, 
    64.37842, 64.42947, 64.45742, 64.46261, 64.44549, 64.40664, 64.34672, 
    64.26649, 64.16679, 64.04854, 63.91275, 63.76048, 63.59284, 63.41101, 
    63.21621, 63.00968, 62.79271, 62.56661, 62.33272, 62.09239, 61.84698, 
    61.5979, 61.34653, 61.09428, 60.84259, 60.59286, 60.34655, 60.10511, 
    59.86998, 59.64262, 59.42447, 59.21699, 59.02159, 58.83967, 58.67258, 
    58.52162, 58.38801, 58.27287, 58.17719, 58.10183, 58.0475, 58.01469, 
    58.00372, 58.01469, 58.0475, 58.10183, 58.17719, 58.27287, 58.38801, 
    58.52162, 58.67258, 58.83967, 59.02159, 59.21699, 59.42447, 59.64262, 
    59.86998, 60.10511, 60.34655, 60.59286, 60.84259, 61.09428, 61.34653, 
    61.5979, 61.84698, 62.09239, 62.33272, 62.56661, 62.79271, 63.00968, 
    63.21621, 63.41101, 63.59284, 63.76048, 63.91275, 64.04854, 64.16679, 
    64.26649, 64.34672, 64.40664, 64.44549, 64.46261, 64.45742, 64.42947, 
    64.37842, 64.304, 64.20609, 64.08468, 63.93984, 63.77176, 63.58075, 
    63.3672, 63.13157, 62.87445, 62.59647, 62.29833, 61.98082, 61.64475, 
    61.291, 60.9205, 60.53419, 60.13306, 59.71813, 59.29044, 58.85105, 
    58.40106, 57.94158, 57.47375, 56.99876, 56.51779, 56.03211, 55.54301, 
    55.05185, 54.56006, 54.06915, 53.58073, 53.09655, 52.61848, 52.14857, 
    51.68906, 51.2424, 50.8113, 50.39874, 50.00798, 49.64257, 49.3063, 
    49.00319, 48.73734, 48.51285, 48.33353, 48.20277, 48.12318, 48.09645,
  48.32068, 48.29103, 48.32068, 48.40891, 48.55354, 48.75123, 48.9978, 
    49.28855, 49.61863, 49.98325, 50.37781, 50.7981, 51.24025, 51.70077, 
    52.17654, 52.66476, 53.16291, 53.66874, 54.18018, 54.69537, 55.21259, 
    55.73024, 56.24681, 56.76091, 57.27117, 57.77631, 58.27507, 58.76625, 
    59.24865, 59.72111, 60.18249, 60.63166, 61.06752, 61.48898, 61.89495, 
    62.2844, 62.65631, 63.00969, 63.34359, 63.65711, 63.94939, 64.21967, 
    64.4672, 64.69138, 64.89165, 65.06756, 65.21877, 65.34507, 65.44633, 
    65.52256, 65.57391, 65.60062, 65.60308, 65.58179, 65.53739, 65.47059, 
    65.38222, 65.27322, 65.14459, 64.99744, 64.83292, 64.65224, 64.45668, 
    64.24754, 64.02619, 63.79399, 63.55234, 63.30267, 63.04639, 62.78497, 
    62.51986, 62.25252, 61.98443, 61.71707, 61.45193, 61.19053, 60.93434, 
    60.6849, 60.44372, 60.21231, 59.99218, 59.78484, 59.59175, 59.41435, 
    59.25401, 59.11205, 58.98967, 58.88793, 58.80779, 58.74997, 58.71506, 
    58.70338, 58.71506, 58.74997, 58.80779, 58.88793, 58.98967, 59.11205, 
    59.25401, 59.41435, 59.59175, 59.78484, 59.99218, 60.21231, 60.44372, 
    60.6849, 60.93434, 61.19053, 61.45193, 61.71707, 61.98443, 62.25252, 
    62.51986, 62.78497, 63.04639, 63.30267, 63.55234, 63.79399, 64.02619, 
    64.24754, 64.45668, 64.65224, 64.83292, 64.99744, 65.14459, 65.27322, 
    65.38222, 65.47059, 65.53739, 65.58179, 65.60308, 65.60062, 65.57391, 
    65.52256, 65.44633, 65.34507, 65.21877, 65.06756, 64.89165, 64.69138, 
    64.4672, 64.21967, 63.94939, 63.65711, 63.34359, 63.00969, 62.65631, 
    62.2844, 61.89495, 61.48898, 61.06752, 60.63166, 60.18249, 59.72111, 
    59.24865, 58.76625, 58.27507, 57.77631, 57.27117, 56.76091, 56.24681, 
    55.73024, 55.21259, 54.69537, 54.18018, 53.66874, 53.16291, 52.66476, 
    52.17654, 51.70077, 51.24025, 50.7981, 50.37781, 49.98325, 49.61863, 
    49.28855, 48.9978, 48.75123, 48.55354, 48.40891, 48.32068, 48.29103,
  48.49963, 48.46671, 48.49963, 48.59744, 48.75734, 48.97508, 49.24543, 
    49.5627, 49.9211, 50.31509, 50.73953, 51.18976, 51.66163, 52.15149, 
    52.65608, 53.17257, 53.69843, 54.23139, 54.76944, 55.31073, 55.85358, 
    56.39642, 56.93778, 57.47627, 58.01056, 58.53938, 59.06146, 59.57561, 
    60.08062, 60.5753, 61.0585, 61.52904, 61.98578, 62.42758, 62.8533, 
    63.26183, 63.65208, 64.02298, 64.37351, 64.70267, 65.00952, 65.29321, 
    65.55291, 65.78793, 65.99763, 66.18151, 66.33916, 66.47034, 66.57487, 
    66.65276, 66.70414, 66.7293, 66.72864, 66.70272, 66.65221, 66.57793, 
    66.48079, 66.36181, 66.22211, 66.06287, 65.88538, 65.69096, 65.481, 
    65.25689, 65.0201, 64.77209, 64.51437, 64.24844, 63.97581, 63.69802, 
    63.41657, 63.13302, 62.84889, 62.56573, 62.28509, 62.00851, 61.73756, 
    61.47382, 61.21884, 60.97421, 60.74149, 60.52226, 60.31806, 60.1304, 
    59.96074, 59.81046, 59.68086, 59.57309, 59.48816, 59.42689, 59.38988, 
    59.3775, 59.38988, 59.42689, 59.48816, 59.57309, 59.68086, 59.81046, 
    59.96074, 60.1304, 60.31806, 60.52226, 60.74149, 60.97421, 61.21884, 
    61.47382, 61.73756, 62.00851, 62.28509, 62.56573, 62.84889, 63.13302, 
    63.41657, 63.69802, 63.97581, 64.24844, 64.51437, 64.77209, 65.0201, 
    65.25689, 65.481, 65.69096, 65.88538, 66.06287, 66.22211, 66.36181, 
    66.48079, 66.57793, 66.65221, 66.70272, 66.72864, 66.7293, 66.70414, 
    66.65276, 66.57487, 66.47034, 66.33916, 66.18151, 65.99763, 65.78793, 
    65.55291, 65.29321, 65.00952, 64.70267, 64.37351, 64.02298, 63.65208, 
    63.26183, 62.8533, 62.42758, 61.98578, 61.52904, 61.0585, 60.5753, 
    60.08062, 59.57561, 59.06146, 58.53938, 58.01056, 57.47627, 56.93778, 
    56.39642, 55.85358, 55.31073, 54.76944, 54.23139, 53.69843, 53.17257, 
    52.65608, 52.15149, 51.66163, 51.18976, 50.73953, 50.31509, 49.9211, 
    49.5627, 49.24543, 48.97508, 48.75734, 48.59744, 48.49963, 48.46671,
  48.66188, 48.62529, 48.66188, 48.77037, 48.94714, 49.18674, 49.48269, 
    49.82803, 50.216, 50.64024, 51.09504, 51.57537, 52.07685, 52.59568, 
    53.12859, 53.67271, 54.22554, 54.78488, 55.34874, 55.91534, 56.48304, 
    57.05032, 57.61575, 58.17798, 58.73571, 59.28766, 59.83261, 60.36934, 
    60.89664, 61.41331, 61.91816, 62.40998, 62.88759, 63.34979, 63.79538, 
    64.22318, 64.63201, 65.02072, 65.3882, 65.73335, 66.05512, 66.35257, 
    66.62477, 66.87093, 67.09032, 67.28237, 67.44659, 67.58268, 67.69044, 
    67.76985, 67.82104, 67.84431, 67.84011, 67.80904, 67.75185, 67.66944, 
    67.56281, 67.43311, 67.28156, 67.10947, 66.91824, 66.70931, 66.48419, 
    66.24441, 65.99152, 65.72712, 65.45279, 65.17012, 64.88072, 64.58619, 
    64.28812, 63.98813, 63.68779, 63.38871, 63.0925, 62.80074, 62.51506, 
    62.23706, 61.96837, 61.71062, 61.46544, 61.23445, 61.01926, 60.82146, 
    60.64257, 60.48408, 60.34735, 60.23361, 60.14395, 60.07924, 60.04015, 
    60.02708, 60.04015, 60.07924, 60.14395, 60.23361, 60.34735, 60.48408, 
    60.64257, 60.82146, 61.01926, 61.23445, 61.46544, 61.71062, 61.96837, 
    62.23706, 62.51506, 62.80074, 63.0925, 63.38871, 63.68779, 63.98813, 
    64.28812, 64.58619, 64.88072, 65.17012, 65.45279, 65.72712, 65.99152, 
    66.24441, 66.48419, 66.70931, 66.91824, 67.10947, 67.28156, 67.43311, 
    67.56281, 67.66944, 67.75185, 67.80904, 67.84011, 67.84431, 67.82104, 
    67.76985, 67.69044, 67.58268, 67.44659, 67.28237, 67.09032, 66.87093, 
    66.62477, 66.35257, 66.05512, 65.73335, 65.3882, 65.02072, 64.63201, 
    64.22318, 63.79538, 63.34979, 62.88759, 62.40998, 61.91816, 61.41331, 
    60.89664, 60.36934, 59.83261, 59.28766, 58.73571, 58.17798, 57.61575, 
    57.05032, 56.48304, 55.91534, 55.34874, 54.78488, 54.22554, 53.67271, 
    53.12859, 52.59568, 52.07685, 51.57537, 51.09504, 50.64024, 50.216, 
    49.82803, 49.48269, 49.18674, 48.94714, 48.77037, 48.66188, 48.62529,
  48.80913, 48.76841, 48.80913, 48.92957, 49.125, 49.38846, 49.71184, 
    50.08679, 50.50539, 50.96051, 51.44589, 51.9562, 52.48689, 53.0341, 
    53.59457, 54.16548, 54.7444, 55.32918, 55.91793, 56.50894, 57.10062, 
    57.69153, 58.28027, 58.86554, 59.44607, 60.02061, 60.58795, 61.14686, 
    61.69614, 62.23457, 62.76093, 63.27398, 63.77248, 64.25519, 64.72083, 
    65.16814, 65.59587, 66.00276, 66.38759, 66.74916, 67.08632, 67.39797, 
    67.68311, 67.9408, 68.17024, 68.37073, 68.54173, 68.68282, 68.79381, 
    68.87462, 68.92539, 68.94643, 68.93822, 68.90145, 68.83694, 68.74567, 
    68.62879, 68.48755, 68.3233, 68.13749, 67.93166, 67.70741, 67.46633, 
    67.21012, 66.94045, 66.65901, 66.36749, 66.06759, 65.76099, 65.44938, 
    65.13441, 64.81776, 64.50108, 64.18601, 63.8742, 63.5673, 63.26696, 
    62.97483, 62.69258, 62.42189, 62.16443, 61.92188, 61.6959, 61.48815, 
    61.30023, 61.13368, 60.98996, 60.87037, 60.77607, 60.70799, 60.66686, 
    60.6531, 60.66686, 60.70799, 60.77607, 60.87037, 60.98996, 61.13368, 
    61.30023, 61.48815, 61.6959, 61.92188, 62.16443, 62.42189, 62.69258, 
    62.97483, 63.26696, 63.5673, 63.8742, 64.18601, 64.50108, 64.81776, 
    65.13441, 65.44938, 65.76099, 66.06759, 66.36749, 66.65901, 66.94045, 
    67.21012, 67.46633, 67.70741, 67.93166, 68.13749, 68.3233, 68.48755, 
    68.62879, 68.74567, 68.83694, 68.90145, 68.93822, 68.94643, 68.92539, 
    68.87462, 68.79381, 68.68282, 68.54173, 68.37073, 68.17024, 67.9408, 
    67.68311, 67.39797, 67.08632, 66.74916, 66.38759, 66.00276, 65.59587, 
    65.16814, 64.72083, 64.25519, 63.77248, 63.27398, 62.76093, 62.23457, 
    61.69614, 61.14686, 60.58795, 60.02061, 59.44607, 58.86554, 58.28027, 
    57.69153, 57.10062, 56.50894, 55.91793, 55.32918, 54.7444, 54.16548, 
    53.59457, 53.0341, 52.48689, 51.9562, 51.44589, 50.96051, 50.50539, 
    50.08679, 49.71184, 49.38846, 49.125, 48.92957, 48.80913, 48.76841,
  48.94296, 48.89758, 48.94296, 49.07684, 49.29296, 49.58239, 49.93505, 
    50.34097, 50.79105, 51.27737, 51.79324, 52.33308, 52.89229, 53.46704, 
    54.0541, 54.65078, 55.25472, 55.86391, 56.47653, 57.09095, 57.70569, 
    58.31934, 58.9306, 59.53818, 60.14086, 60.73742, 61.32665, 61.90735, 
    62.4783, 63.03828, 63.58602, 64.12027, 64.63973, 65.1431, 65.62903, 
    66.09618, 66.54319, 66.96871, 67.37141, 67.74994, 68.10303, 68.42947, 
    68.72808, 68.99783, 69.23775, 69.44706, 69.62509, 69.77138, 69.88563, 
    69.96776, 70.01788, 70.03633, 70.02364, 69.98056, 69.90802, 69.80711, 
    69.67911, 69.5254, 69.34751, 69.14704, 68.92569, 68.68518, 68.4273, 
    68.15385, 67.86665, 67.56749, 67.25819, 66.94055, 66.61633, 66.28728, 
    65.95516, 65.62167, 65.28853, 64.95743, 64.63006, 64.3081, 63.99323, 
    63.68716, 63.39157, 63.10819, 62.83872, 62.58489, 62.34842, 62.131, 
    61.9343, 61.75994, 61.60944, 61.48418, 61.38538, 61.31404, 61.27094, 
    61.25651, 61.27094, 61.31404, 61.38538, 61.48418, 61.60944, 61.75994, 
    61.9343, 62.131, 62.34842, 62.58489, 62.83872, 63.10819, 63.39157, 
    63.68716, 63.99323, 64.3081, 64.63006, 64.95743, 65.28853, 65.62167, 
    65.95516, 66.28728, 66.61633, 66.94055, 67.25819, 67.56749, 67.86665, 
    68.15385, 68.4273, 68.68518, 68.92569, 69.14704, 69.34751, 69.5254, 
    69.67911, 69.80711, 69.90802, 69.98056, 70.02364, 70.03633, 70.01788, 
    69.96776, 69.88563, 69.77138, 69.62509, 69.44706, 69.23775, 68.99783, 
    68.72808, 68.42947, 68.10303, 67.74994, 67.37141, 66.96871, 66.54319, 
    66.09618, 65.62903, 65.1431, 64.63973, 64.12027, 63.58602, 63.03828, 
    62.4783, 61.90735, 61.32665, 60.73742, 60.14086, 59.53818, 58.9306, 
    58.31934, 57.70569, 57.09095, 56.47653, 55.86391, 55.25472, 54.65078, 
    54.0541, 53.46704, 52.89229, 52.33308, 51.79324, 51.27737, 50.79105, 
    50.34097, 49.93505, 49.58239, 49.29296, 49.07684, 48.94296, 48.89758,
  49.06485, 49.01415, 49.06485, 49.21389, 49.45297, 49.77058, 50.1543, 
    50.59235, 51.07442, 51.59192, 52.13781, 52.70642, 53.29319, 53.89436, 
    54.50686, 55.1281, 55.75589, 56.38832, 57.0237, 57.66049, 58.29729, 
    58.93279, 59.56571, 60.19484, 60.819, 61.43699, 62.04763, 62.64973, 
    63.24205, 63.82336, 64.3924, 64.94785, 65.48837, 66.01259, 66.5191, 
    67.00648, 67.47325, 67.91795, 68.33912, 68.73528, 69.10499, 69.44689, 
    69.75967, 70.04209, 70.29308, 70.5117, 70.69714, 70.84886, 70.96648, 
    71.04987, 71.09912, 71.11461, 71.09691, 71.04685, 70.96549, 70.85405, 
    70.71396, 70.54678, 70.35421, 70.13803, 69.90012, 69.64237, 69.36674, 
    69.07519, 68.76965, 68.45208, 68.12439, 67.78848, 67.44621, 67.0994, 
    66.74987, 66.39939, 66.04972, 65.7026, 65.35974, 65.02287, 64.69369, 
    64.37392, 64.0653, 63.76956, 63.48844, 63.22371, 62.97711, 62.7504, 
    62.54529, 62.36346, 62.20647, 62.07579, 61.9727, 61.89826, 61.85326, 
    61.83821, 61.85326, 61.89826, 61.9727, 62.07579, 62.20647, 62.36346, 
    62.54529, 62.7504, 62.97711, 63.22371, 63.48844, 63.76956, 64.0653, 
    64.37392, 64.69369, 65.02287, 65.35974, 65.7026, 66.04972, 66.39939, 
    66.74987, 67.0994, 67.44621, 67.78848, 68.12439, 68.45208, 68.76965, 
    69.07519, 69.36674, 69.64237, 69.90012, 70.13803, 70.35421, 70.54678, 
    70.71396, 70.85405, 70.96549, 71.04685, 71.09691, 71.11461, 71.09912, 
    71.04987, 70.96648, 70.84886, 70.69714, 70.5117, 70.29308, 70.04209, 
    69.75967, 69.44689, 69.10499, 68.73528, 68.33912, 67.91795, 67.47325, 
    67.00648, 66.5191, 66.01259, 65.48837, 64.94785, 64.3924, 63.82336, 
    63.24205, 62.64973, 62.04763, 61.43699, 60.819, 60.19484, 59.56571, 
    58.93279, 58.29729, 57.66049, 57.0237, 56.38832, 55.75589, 55.1281, 
    54.50686, 53.89436, 53.29319, 52.70642, 52.13781, 51.59192, 51.07442, 
    50.59235, 50.1543, 49.77058, 49.45297, 49.21389, 49.06485, 49.01415,
  49.17618, 49.11938, 49.17618, 49.34239, 49.60692, 49.95499, 50.37137, 
    50.84236, 51.35654, 51.90476, 52.47985, 53.07615, 53.68922, 54.31551, 
    54.95209, 55.59658, 56.24692, 56.90136, 57.55832, 58.21637, 58.87421, 
    59.53059, 60.18432, 60.83424, 61.47919, 62.11802, 62.74957, 63.37265, 
    63.98605, 64.58852, 65.17875, 65.75542, 66.31713, 66.86246, 67.38992, 
    67.89796, 68.38506, 68.84958, 69.28993, 69.70449, 70.09165, 70.44985, 
    70.77761, 71.07351, 71.33628, 71.56481, 71.75816, 71.91565, 72.0368, 
    72.12142, 72.16961, 72.18173, 72.15844, 72.10067, 72.0096, 71.88663, 
    71.73337, 71.55157, 71.34315, 71.11011, 70.8545, 70.57844, 70.28404, 
    69.97344, 69.64874, 69.31202, 68.96531, 68.6106, 68.24986, 67.88498, 
    67.51783, 67.15025, 66.78403, 66.42094, 66.06273, 65.71115, 65.36793, 
    65.03481, 64.71353, 64.40585, 64.11353, 63.83837, 63.58213, 63.34661, 
    63.13356, 62.94469, 62.78163, 62.64589, 62.53879, 62.46144, 62.41469, 
    62.39905, 62.41469, 62.46144, 62.53879, 62.64589, 62.78163, 62.94469, 
    63.13356, 63.34661, 63.58213, 63.83837, 64.11353, 64.40585, 64.71353, 
    65.03481, 65.36793, 65.71115, 66.06273, 66.42094, 66.78403, 67.15025, 
    67.51783, 67.88498, 68.24986, 68.6106, 68.96531, 69.31202, 69.64874, 
    69.97344, 70.28404, 70.57844, 70.8545, 71.11011, 71.34315, 71.55157, 
    71.73337, 71.88663, 72.0096, 72.10067, 72.15844, 72.18173, 72.16961, 
    72.12142, 72.0368, 71.91565, 71.75816, 71.56481, 71.33628, 71.07351, 
    70.77761, 70.44985, 70.09165, 69.70449, 69.28993, 68.84958, 68.38506, 
    67.89796, 67.38992, 66.86246, 66.31713, 65.75542, 65.17875, 64.58852, 
    63.98605, 63.37265, 62.74957, 62.11802, 61.47919, 60.83424, 60.18432, 
    59.53059, 58.87421, 58.21637, 57.55832, 56.90136, 56.24692, 55.59658, 
    54.95209, 54.31551, 53.68922, 53.07615, 52.47985, 51.90476, 51.35654, 
    50.84236, 50.37137, 49.95499, 49.60692, 49.34239, 49.17618, 49.11938,
  49.27823, 49.21439, 49.27823, 49.46397, 49.75667, 50.1374, 50.58774, 
    51.09206, 51.63798, 52.21606, 52.81913, 53.44172, 54.07962, 54.7295, 
    55.38869, 56.05498, 56.72651, 57.40165, 58.07897, 58.75715, 59.43497, 
    60.11127, 60.78493, 61.45483, 62.11987, 62.77893, 63.43088, 64.07455, 
    64.70872, 65.33213, 65.94349, 66.54141, 67.12448, 67.69118, 68.23998, 
    68.76924, 69.27728, 69.76237, 70.22274, 70.65661, 71.06217, 71.43768, 
    71.7814, 72.09173, 72.36716, 72.60638, 72.80828, 72.97198, 73.09691, 
    73.18279, 73.22971, 73.23804, 73.20851, 73.14219, 73.04041, 72.90478, 
    72.73711, 72.53943, 72.31386, 72.06265, 71.7881, 71.49254, 71.17829, 
    70.84766, 70.50291, 70.14628, 69.7799, 69.40588, 69.02627, 68.64303, 
    68.25809, 67.87333, 67.49058, 67.11164, 66.73829, 66.37228, 66.01537, 
    65.6693, 65.33584, 65.01673, 64.71378, 64.42876, 64.16349, 63.91976, 
    63.69936, 63.50402, 63.3354, 63.19505, 63.08432, 63.00436, 62.95603, 
    62.93986, 62.95603, 63.00436, 63.08432, 63.19505, 63.3354, 63.50402, 
    63.69936, 63.91976, 64.16349, 64.42876, 64.71378, 65.01673, 65.33584, 
    65.6693, 66.01537, 66.37228, 66.73829, 67.11164, 67.49058, 67.87333, 
    68.25809, 68.64303, 69.02627, 69.40588, 69.7799, 70.14628, 70.50291, 
    70.84766, 71.17829, 71.49254, 71.7881, 72.06265, 72.31386, 72.53943, 
    72.73711, 72.90478, 73.04041, 73.14219, 73.20851, 73.23804, 73.22971, 
    73.18279, 73.09691, 72.97198, 72.80828, 72.60638, 72.36716, 72.09173, 
    71.7814, 71.43768, 71.06217, 70.65661, 70.22274, 69.76237, 69.27728, 
    68.76924, 68.23998, 67.69118, 67.12448, 66.54141, 65.94349, 65.33213, 
    64.70872, 64.07455, 63.43088, 62.77893, 62.11987, 61.45483, 60.78493, 
    60.11127, 59.43497, 58.75715, 58.07897, 57.40165, 56.72651, 56.05498, 
    55.38869, 54.7295, 54.07962, 53.44172, 52.81913, 52.21606, 51.63798, 
    51.09206, 50.58774, 50.1374, 49.75667, 49.46397, 49.27823, 49.21439,
  49.37224, 49.30021, 49.37224, 49.58023, 49.904, 50.31941, 50.80456, 
    51.34202, 51.91881, 52.52541, 53.1549, 53.80212, 54.46316, 55.13499, 
    55.8152, 56.50179, 57.19306, 57.88757, 58.584, 59.28114, 59.97787, 
    60.67311, 61.36579, 62.05486, 62.73927, 63.41795, 64.08977, 64.75359, 
    65.40821, 66.05238, 66.68476, 67.30399, 67.90856, 68.49696, 69.06752, 
    69.61855, 70.14825, 70.65473, 71.13608, 71.5903, 72.0154, 72.40937, 
    72.77025, 73.09615, 73.38533, 73.6362, 73.84741, 74.01791, 74.14697, 
    74.2342, 74.27963, 74.28371, 74.24722, 74.17139, 74.05777, 73.90817, 
    73.72472, 73.50969, 73.26551, 72.99471, 72.69984, 72.3835, 72.04823, 
    71.69652, 71.33082, 70.95349, 70.56682, 70.17299, 69.77414, 69.3723, 
    68.96944, 68.56749, 68.1683, 67.7737, 67.38547, 67.00539, 66.63522, 
    66.2767, 65.9316, 65.60169, 65.28876, 64.99459, 64.721, 64.4698, 
    64.24277, 64.04167, 63.86816, 63.72379, 63.60992, 63.52772, 63.47803, 
    63.46141, 63.47803, 63.52772, 63.60992, 63.72379, 63.86816, 64.04167, 
    64.24277, 64.4698, 64.721, 64.99459, 65.28876, 65.60169, 65.9316, 
    66.2767, 66.63522, 67.00539, 67.38547, 67.7737, 68.1683, 68.56749, 
    68.96944, 69.3723, 69.77414, 70.17299, 70.56682, 70.95349, 71.33082, 
    71.69652, 72.04823, 72.3835, 72.69984, 72.99471, 73.26551, 73.50969, 
    73.72472, 73.90817, 74.05777, 74.17139, 74.24722, 74.28371, 74.27963, 
    74.2342, 74.14697, 74.01791, 73.84741, 73.6362, 73.38533, 73.09615, 
    72.77025, 72.40937, 72.0154, 71.5903, 71.13608, 70.65473, 70.14825, 
    69.61855, 69.06752, 68.49696, 67.90856, 67.30399, 66.68476, 66.05238, 
    65.40821, 64.75359, 64.08977, 63.41795, 62.73927, 62.05486, 61.36579, 
    60.67311, 59.97787, 59.28114, 58.584, 57.88757, 57.19306, 56.50179, 
    55.8152, 55.13499, 54.46316, 53.80212, 53.1549, 52.52541, 51.91881, 
    51.34202, 50.80456, 50.31941, 49.904, 49.58023, 49.37224, 49.30021,
  49.45941, 49.37779, 49.45941, 49.6928, 50.05057, 50.5023, 51.02249, 
    51.59231, 52.19854, 52.83192, 53.48596, 54.15591, 54.83826, 55.5303, 
    56.22986, 56.93518, 57.64476, 58.35727, 59.07154, 59.78647, 60.50102, 
    61.21419, 61.92498, 62.6324, 63.33544, 64.03307, 64.72421, 65.40772, 
    66.08245, 66.74713, 67.40044, 68.04098, 68.66723, 69.2776, 69.8704, 
    70.44381, 70.99592, 71.52472, 72.02809, 72.50386, 72.94978, 73.36357, 
    73.743, 74.08585, 74.39007, 74.65376, 74.87528, 75.05333, 75.18697, 
    75.27569, 75.31947, 75.31876, 75.27449, 75.18806, 75.06125, 74.89622, 
    74.69537, 74.46134, 74.19691, 73.90493, 73.58826, 73.24976, 72.89221, 
    72.51835, 72.13076, 71.73198, 71.32439, 70.91029, 70.49188, 70.07125, 
    69.65042, 69.23133, 68.81586, 68.40585, 68.00311, 67.60939, 67.22646, 
    66.85609, 66.50001, 66.16, 65.83785, 65.53535, 65.2543, 64.99651, 
    64.76374, 64.55775, 64.38016, 64.23251, 64.11614, 64.03217, 63.98144, 
    63.96447, 63.98144, 64.03217, 64.11614, 64.23251, 64.38016, 64.55775, 
    64.76374, 64.99651, 65.2543, 65.53535, 65.83785, 66.16, 66.50001, 
    66.85609, 67.22646, 67.60939, 68.00311, 68.40585, 68.81586, 69.23133, 
    69.65042, 70.07125, 70.49188, 70.91029, 71.32439, 71.73198, 72.13076, 
    72.51835, 72.89221, 73.24976, 73.58826, 73.90493, 74.19691, 74.46134, 
    74.69537, 74.89622, 75.06125, 75.18806, 75.27449, 75.31876, 75.31947, 
    75.27569, 75.18697, 75.05333, 74.87528, 74.65376, 74.39007, 74.08585, 
    73.743, 73.36357, 72.94978, 72.50386, 72.02809, 71.52472, 70.99592, 
    70.44381, 69.8704, 69.2776, 68.66723, 68.04098, 67.40044, 66.74713, 
    66.08245, 65.40772, 64.72421, 64.03307, 63.33544, 62.6324, 61.92498, 
    61.21419, 60.50102, 59.78647, 59.07154, 58.35727, 57.64476, 56.93518, 
    56.22986, 55.5303, 54.83826, 54.15591, 53.48596, 52.83192, 52.19854, 
    51.59231, 51.02249, 50.5023, 50.05057, 49.6928, 49.45941, 49.37779,
  49.54091, 49.44797, 49.54091, 49.80328, 50.19788, 50.68695, 51.24167, 
    51.84238, 52.4761, 53.13417, 53.81063, 54.50129, 55.20302, 55.91344, 
    56.63068, 57.35317, 58.07958, 58.80874, 59.53959, 60.27112, 61.00239, 
    61.73247, 62.46043, 63.18534, 63.90624, 64.62214, 65.33199, 66.03472, 
    66.72916, 67.41407, 68.08815, 68.74997, 69.39802, 70.03065, 70.64612, 
    71.24252, 71.81785, 72.36993, 72.89648, 73.3951, 73.8633, 74.29848, 
    74.69807, 75.05951, 75.38034, 75.65829, 75.89136, 76.0779, 76.21672, 
    76.30715, 76.34908, 76.34301, 76.29001, 76.19169, 76.05016, 75.86795, 
    75.64788, 75.393, 75.10648, 74.79156, 74.45145, 74.08932, 73.70821, 
    73.31107, 72.90068, 72.47969, 72.05063, 71.61586, 71.17764, 70.73811, 
    70.29932, 69.86323, 69.43173, 69.00666, 68.58983, 68.183, 67.78792, 
    67.40635, 67.04004, 66.69075, 66.36026, 66.05036, 65.76284, 65.49947, 
    65.26202, 65.05217, 64.87152, 64.72152, 64.60344, 64.51832, 64.46693, 
    64.44975, 64.46693, 64.51832, 64.60344, 64.72152, 64.87152, 65.05217, 
    65.26202, 65.49947, 65.76284, 66.05036, 66.36026, 66.69075, 67.04004, 
    67.40635, 67.78792, 68.183, 68.58983, 69.00666, 69.43173, 69.86323, 
    70.29932, 70.73811, 71.17764, 71.61586, 72.05063, 72.47969, 72.90068, 
    73.31107, 73.70821, 74.08932, 74.45145, 74.79156, 75.10648, 75.393, 
    75.64788, 75.86795, 76.05016, 76.19169, 76.29001, 76.34301, 76.34908, 
    76.30715, 76.21672, 76.0779, 75.89136, 75.65829, 75.38034, 75.05951, 
    74.69807, 74.29848, 73.8633, 73.3951, 72.89648, 72.36993, 71.81785, 
    71.24252, 70.64612, 70.03065, 69.39802, 68.74997, 68.08815, 67.41407, 
    66.72916, 66.03472, 65.33199, 64.62214, 63.90624, 63.18534, 62.46043, 
    61.73247, 61.00239, 60.27112, 59.53959, 58.80874, 58.07958, 57.35317, 
    56.63068, 55.91344, 55.20302, 54.50129, 53.81063, 53.13417, 52.4761, 
    51.84238, 51.24167, 50.68695, 50.19788, 49.80328, 49.54091, 49.44797,
  49.61793, 49.51152, 49.61793, 49.91324, 50.34711, 50.8737, 51.46157, 
    52.09106, 52.74991, 53.43027, 54.1269, 54.83612, 55.55526, 56.28226, 
    57.01549, 57.75359, 58.49538, 59.23983, 59.98599, 60.73295, 61.47984, 
    62.2258, 62.96998, 63.71149, 64.44943, 65.18286, 65.91079, 66.63216, 
    67.34585, 68.05064, 68.74525, 69.42828, 70.09817, 70.75328, 71.39182, 
    72.01181, 72.61115, 73.18752, 73.73848, 74.26139, 74.75346, 75.21181, 
    75.63345, 76.0154, 76.35472, 76.64868, 76.89481, 77.09103, 77.23584, 
    77.3283, 77.36822, 77.3561, 77.29323, 77.1815, 77.02345, 76.82204, 
    76.58063, 76.30276, 75.9921, 75.65231, 75.28703, 74.89972, 74.49372, 
    74.0722, 73.63811, 73.19424, 72.7432, 72.28745, 71.82926, 71.37083, 
    70.91421, 70.46135, 70.01417, 69.57448, 69.14408, 68.72473, 68.31819, 
    67.92619, 67.55048, 67.19282, 66.85497, 66.53873, 66.24585, 65.9781, 
    65.73719, 65.52473, 65.34222, 65.191, 65.0722, 64.98671, 64.93516, 
    64.91794, 64.93516, 64.98671, 65.0722, 65.191, 65.34222, 65.52473, 
    65.73719, 65.9781, 66.24585, 66.53873, 66.85497, 67.19282, 67.55048, 
    67.92619, 68.31819, 68.72473, 69.14408, 69.57448, 70.01417, 70.46135, 
    70.91421, 71.37083, 71.82926, 72.28745, 72.7432, 73.19424, 73.63811, 
    74.0722, 74.49372, 74.89972, 75.28703, 75.65231, 75.9921, 76.30276, 
    76.58063, 76.82204, 77.02345, 77.1815, 77.29323, 77.3561, 77.36822, 
    77.3283, 77.23584, 77.09103, 76.89481, 76.64868, 76.35472, 76.0154, 
    75.63345, 75.21181, 74.75346, 74.26139, 73.73848, 73.18752, 72.61115, 
    72.01181, 71.39182, 70.75328, 70.09817, 69.42828, 68.74525, 68.05064, 
    67.34585, 66.63216, 65.91079, 65.18286, 64.44943, 63.71149, 62.96998, 
    62.2258, 61.47984, 60.73295, 59.98599, 59.23983, 58.49538, 57.75359, 
    57.01549, 56.28226, 55.55526, 54.83612, 54.1269, 53.43027, 52.74991, 
    52.09106, 51.46157, 50.8737, 50.34711, 49.91324, 49.61793, 49.51152,
  49.6917, 49.56914, 49.6917, 50.02419, 50.499, 51.06221, 51.68102, 52.33659, 
    53.01786, 53.71797, 54.43241, 55.15807, 55.89267, 56.63445, 57.38202, 
    58.1342, 58.88995, 59.64837, 60.40858, 61.16979, 61.93119, 62.69198, 
    63.45139, 64.20857, 64.9627, 65.71288, 66.45815, 67.19753, 67.92991, 
    68.65414, 69.36897, 70.07298, 70.76467, 71.44238, 72.10429, 72.74841, 
    73.3725, 73.97417, 74.55079, 75.0995, 75.61723, 76.10072, 76.54655, 
    76.95124, 77.3113, 77.62341, 77.88448, 78.09192, 78.24372, 78.33866, 
    78.37637, 78.35744, 78.28333, 78.15639, 77.97964, 77.75668, 77.49148, 
    77.18821, 76.85112, 76.48439, 76.09206, 75.67799, 75.24577, 74.79881, 
    74.34021, 73.87288, 73.39951, 72.92257, 72.4444, 71.96718, 71.49297, 
    71.0237, 70.56128, 70.10751, 69.66416, 69.233, 68.81575, 68.41416, 
    68.02996, 67.66492, 67.3208, 66.99937, 66.7024, 66.4316, 66.18863, 
    65.97501, 65.79209, 65.64104, 65.52274, 65.43783, 65.38674, 65.36969, 
    65.38674, 65.43783, 65.52274, 65.64104, 65.79209, 65.97501, 66.18863, 
    66.4316, 66.7024, 66.99937, 67.3208, 67.66492, 68.02996, 68.41416, 
    68.81575, 69.233, 69.66416, 70.10751, 70.56128, 71.0237, 71.49297, 
    71.96718, 72.4444, 72.92257, 73.39951, 73.87288, 74.34021, 74.79881, 
    75.24577, 75.67799, 76.09206, 76.48439, 76.85112, 77.18821, 77.49148, 
    77.75668, 77.97964, 78.15639, 78.28333, 78.35744, 78.37637, 78.33866, 
    78.24372, 78.09192, 77.88448, 77.62341, 77.3113, 76.95124, 76.54655, 
    76.10072, 75.61723, 75.0995, 74.55079, 73.97417, 73.3725, 72.74841, 
    72.10429, 71.44238, 70.76467, 70.07298, 69.36897, 68.65414, 67.92991, 
    67.19753, 66.45815, 65.71288, 64.9627, 64.20857, 63.45139, 62.69198, 
    61.93119, 61.16979, 60.40858, 59.64837, 58.88995, 58.1342, 57.38202, 
    56.63445, 55.89267, 55.15807, 54.43241, 53.71797, 53.01786, 52.33659, 
    51.68102, 51.06221, 50.499, 50.02419, 49.6917, 49.56914,
  49.7635, 49.62147, 49.7635, 50.13739, 50.65365, 51.2514, 51.89813, 52.5767, 
    53.27751, 53.99475, 54.72467, 55.46467, 56.21283, 56.96767, 57.728, 
    58.49277, 59.26111, 60.03218, 60.80522, 61.57949, 62.35427, 63.12884, 
    63.90245, 64.67434, 65.44373, 66.20978, 66.9716, 67.72823, 68.47866, 
    69.22176, 69.95632, 70.68099, 71.39429, 72.09459, 72.78005, 73.44867, 
    74.09818, 74.72607, 75.32958, 75.90564, 76.45088, 76.96168, 77.43413, 
    77.86417, 78.24763, 78.58047, 78.85883, 79.07939, 79.23952, 79.33755, 
    79.37289, 79.34618, 79.2592, 79.11483, 78.9168, 78.66949, 78.37767, 
    78.04628, 77.68024, 77.28433, 76.86305, 76.42063, 75.96095, 75.48759, 
    75.00381, 74.5126, 74.01666, 73.51853, 73.02052, 72.52477, 72.03335, 
    71.54816, 71.07108, 70.60387, 70.14829, 69.70609, 69.27898, 68.86871, 
    68.47701, 68.10565, 67.75641, 67.43106, 67.13136, 66.85899, 66.61555, 
    66.40244, 66.22082, 66.07156, 65.95523, 65.87211, 65.82224, 65.80563, 
    65.82224, 65.87211, 65.95523, 66.07156, 66.22082, 66.40244, 66.61555, 
    66.85899, 67.13136, 67.43106, 67.75641, 68.10565, 68.47701, 68.86871, 
    69.27898, 69.70609, 70.14829, 70.60387, 71.07108, 71.54816, 72.03335, 
    72.52477, 73.02052, 73.51853, 74.01666, 74.5126, 75.00381, 75.48759, 
    75.96095, 76.42063, 76.86305, 77.28433, 77.68024, 78.04628, 78.37767, 
    78.66949, 78.9168, 79.11483, 79.2592, 79.34618, 79.37289, 79.33755, 
    79.23952, 79.07939, 78.85883, 78.58047, 78.24763, 77.86417, 77.43413, 
    76.96168, 76.45088, 75.90564, 75.32958, 74.72607, 74.09818, 73.44867, 
    72.78005, 72.09459, 71.39429, 70.68099, 69.95632, 69.22176, 68.47866, 
    67.72823, 66.9716, 66.20978, 65.44373, 64.67434, 63.90245, 63.12884, 
    62.35427, 61.57949, 60.80522, 60.03218, 59.26111, 58.49277, 57.728, 
    56.96767, 56.21283, 55.46467, 54.72467, 53.99475, 53.27751, 52.5767, 
    51.89813, 51.2514, 50.65365, 50.13739, 49.7635, 49.62147,
  49.83468, 49.66908, 49.83468, 50.25368, 50.81035, 51.4394, 52.11046, 
    52.8087, 53.52612, 54.25795, 55.00111, 55.75345, 56.51337, 57.27963, 
    58.05119, 58.82714, 59.60672, 60.38918, 61.17383, 61.96, 62.74704, 
    63.53428, 64.32103, 65.10661, 65.89027, 66.67123, 67.44869, 68.22174, 
    68.98942, 69.75067, 70.50435, 71.24916, 71.98369, 72.70634, 73.41534, 
    74.10866, 74.78405, 75.43895, 76.07047, 76.67538, 77.25005, 77.79045, 
    78.2922, 78.75056, 79.16058, 79.51729, 79.81586, 80.05197, 80.22216, 
    80.3241, 80.3569, 80.32124, 80.21935, 80.05484, 79.83239, 79.55742, 
    79.23571, 78.87315, 78.47546, 78.04803, 77.59591, 77.12365, 76.63539, 
    76.13487, 75.62544, 75.11012, 74.59165, 74.0725, 73.55497, 73.04117, 
    72.53309, 72.03262, 71.54156, 71.06167, 70.59467, 70.14229, 69.70624, 
    69.28825, 68.89008, 68.51352, 68.16036, 67.83242, 67.53146, 67.25915, 
    67.01701, 66.80629, 66.62793, 66.48241, 66.36983, 66.28991, 66.24222, 
    66.22637, 66.24222, 66.28991, 66.36983, 66.48241, 66.62793, 66.80629, 
    67.01701, 67.25915, 67.53146, 67.83242, 68.16036, 68.51352, 68.89008, 
    69.28825, 69.70624, 70.14229, 70.59467, 71.06167, 71.54156, 72.03262, 
    72.53309, 73.04117, 73.55497, 74.0725, 74.59165, 75.11012, 75.62544, 
    76.13487, 76.63539, 77.12365, 77.59591, 78.04803, 78.47546, 78.87315, 
    79.23571, 79.55742, 79.83239, 80.05484, 80.21935, 80.32124, 80.3569, 
    80.3241, 80.22216, 80.05197, 79.81586, 79.51729, 79.16058, 78.75056, 
    78.2922, 77.79045, 77.25005, 76.67538, 76.07047, 75.43895, 74.78405, 
    74.10866, 73.41534, 72.70634, 71.98369, 71.24916, 70.50435, 69.75067, 
    68.98942, 68.22174, 67.44869, 66.67123, 65.89027, 65.10661, 64.32103, 
    63.53428, 62.74704, 61.96, 61.17383, 60.38918, 59.60672, 58.82714, 
    58.05119, 57.27963, 56.51337, 55.75345, 55.00111, 54.25795, 53.52612, 
    52.8087, 52.11046, 51.4394, 50.81035, 50.25368, 49.83468, 49.66908,
  49.90665, 49.71249, 49.90665, 50.37326, 50.96746, 51.62363, 52.31512, 
    53.02969, 53.76089, 54.5049, 55.25919, 56.02202, 56.79203, 57.56816, 
    58.34951, 59.13531, 59.92484, 60.71745, 61.51251, 62.30942, 63.10757, 
    63.90636, 64.70517, 65.50334, 66.30021, 67.09506, 67.88714, 68.67561, 
    69.4596, 70.23812, 71.01009, 71.77432, 72.52946, 73.27401, 74.00623, 
    74.7242, 75.42567, 76.10811, 76.76856, 77.40368, 78.00961, 78.58199, 
    79.1159, 79.60591, 80.04616, 80.43053, 80.75294, 81.00775, 81.19027, 
    81.29724, 81.32732, 81.28123, 81.16186, 80.97382, 80.72313, 80.41657, 
    80.06125, 79.66417, 79.23196, 78.77071, 78.28595, 77.78255, 77.26486, 
    76.7367, 76.20145, 75.66211, 75.12137, 74.58165, 74.04517, 73.51398, 
    72.98997, 72.47501, 71.97081, 71.4791, 71.00158, 70.53994, 70.09589, 
    69.6712, 69.26762, 68.887, 68.53118, 68.20203, 67.90134, 67.63081, 
    67.39191, 67.18574, 67.01289, 66.87337, 66.76661, 66.69159, 66.64718, 
    66.63248, 66.64718, 66.69159, 66.76661, 66.87337, 67.01289, 67.18574, 
    67.39191, 67.63081, 67.90134, 68.20203, 68.53118, 68.887, 69.26762, 
    69.6712, 70.09589, 70.53994, 71.00158, 71.4791, 71.97081, 72.47501, 
    72.98997, 73.51398, 74.04517, 74.58165, 75.12137, 75.66211, 76.20145, 
    76.7367, 77.26486, 77.78255, 78.28595, 78.77071, 79.23196, 79.66417, 
    80.06125, 80.41657, 80.72313, 80.97382, 81.16186, 81.28123, 81.32732, 
    81.29724, 81.19027, 81.00775, 80.75294, 80.43053, 80.04616, 79.60591, 
    79.1159, 78.58199, 78.00961, 77.40368, 76.76856, 76.10811, 75.42567, 
    74.7242, 74.00623, 73.27401, 72.52946, 71.77432, 71.01009, 70.23812, 
    69.4596, 68.67561, 67.88714, 67.09506, 66.30021, 65.50334, 64.70517, 
    63.90636, 63.10757, 62.30942, 61.51251, 60.71745, 59.92484, 59.13531, 
    58.34951, 57.56816, 56.79203, 56.02202, 55.25919, 54.5049, 53.76089, 
    53.02969, 52.31512, 51.62363, 50.96746, 50.37326, 49.90665, 49.71249,
  49.98074, 49.75218, 49.98074, 50.49529, 51.12246, 51.80101, 52.50899, 
    53.23671, 53.97908, 54.73305, 55.49658, 56.26818, 57.04674, 57.83132, 
    58.62113, 59.41548, 60.21373, 61.0153, 61.8196, 62.62609, 63.43421, 
    64.24342, 65.05312, 65.86275, 66.67169, 67.47929, 68.28486, 69.08765, 
    69.88684, 70.68155, 71.47079, 72.25346, 73.02834, 73.79399, 74.54884, 
    75.29102, 76.01842, 76.72855, 77.4185, 78.08486, 78.72369, 79.33031, 
    79.89935, 80.42465, 80.89934, 81.31594, 81.66674, 81.9443, 82.14217, 
    82.25574, 82.2829, 82.22449, 82.08427, 81.86843, 81.5848, 81.24203, 
    80.84888, 80.4137, 79.9441, 79.44688, 78.92797, 78.39249, 77.84489, 
    77.28899, 76.72813, 76.16521, 75.60283, 75.04328, 74.48869, 73.94098, 
    73.402, 72.87347, 72.35711, 71.85455, 71.36748, 70.89755, 70.44652, 
    70.01612, 69.60821, 69.22466, 68.86742, 68.53844, 68.23962, 67.97271, 
    67.73915, 67.53988, 67.3751, 67.24418, 67.14565, 67.07748, 67.03762, 
    67.02453, 67.03762, 67.07748, 67.14565, 67.24418, 67.3751, 67.53988, 
    67.73915, 67.97271, 68.23962, 68.53844, 68.86742, 69.22466, 69.60821, 
    70.01612, 70.44652, 70.89755, 71.36748, 71.85455, 72.35711, 72.87347, 
    73.402, 73.94098, 74.48869, 75.04328, 75.60283, 76.16521, 76.72813, 
    77.28899, 77.84489, 78.39249, 78.92797, 79.44688, 79.9441, 80.4137, 
    80.84888, 81.24203, 81.5848, 81.86843, 82.08427, 82.22449, 82.2829, 
    82.25574, 82.14217, 81.9443, 81.66674, 81.31594, 80.89934, 80.42465, 
    79.89935, 79.33031, 78.72369, 78.08486, 77.4185, 76.72855, 76.01842, 
    75.29102, 74.54884, 73.79399, 73.02834, 72.25346, 71.47079, 70.68155, 
    69.88684, 69.08765, 68.28486, 67.47929, 66.67169, 65.86275, 65.05312, 
    64.24342, 63.43421, 62.62609, 61.8196, 61.0153, 60.21373, 59.41548, 
    58.62113, 57.83132, 57.04674, 56.26818, 55.49658, 54.73305, 53.97908, 
    53.23671, 52.50899, 51.80101, 51.12246, 50.49529, 49.98074, 49.75218,
  50.05792, 49.78856, 50.05792, 50.61779, 51.27207, 51.96816, 52.68894, 
    53.42694, 54.17815, 54.94013, 55.71118, 56.49005, 57.27575, 58.06747, 
    58.86449, 59.66619, 60.472, 61.28136, 62.09375, 62.90866, 63.7256, 
    64.54404, 65.36349, 66.18338, 67.00318, 67.8223, 68.64011, 69.45595, 
    70.26908, 71.07871, 71.88396, 72.68385, 73.47726, 74.26292, 75.03938, 
    75.80494, 76.55762, 77.29511, 78.01461, 78.7128, 79.3857, 80.02852, 
    80.63553, 81.19992, 81.71375, 82.16798, 82.55286, 82.85847, 83.07582, 
    83.19816, 83.22219, 83.1489, 82.98342, 82.73427, 82.41193, 82.02757, 
    81.59199, 81.11507, 80.60542, 80.07044, 79.51636, 78.94839, 78.37096, 
    77.78775, 77.20197, 76.61634, 76.03331, 75.45501, 74.88342, 74.32034, 
    73.76749, 73.22653, 72.69907, 72.18674, 71.69113, 71.21395, 70.75691, 
    70.32183, 69.9106, 69.52522, 69.16776, 68.84031, 68.54496, 68.28358, 
    68.05765, 67.86792, 67.71413, 67.59476, 67.50717, 67.44801, 67.41405, 
    67.40302, 67.41405, 67.44801, 67.50717, 67.59476, 67.71413, 67.86792, 
    68.05765, 68.28358, 68.54496, 68.84031, 69.16776, 69.52522, 69.9106, 
    70.32183, 70.75691, 71.21395, 71.69113, 72.18674, 72.69907, 73.22653, 
    73.76749, 74.32034, 74.88342, 75.45501, 76.03331, 76.61634, 77.20197, 
    77.78775, 78.37096, 78.94839, 79.51636, 80.07044, 80.60542, 81.11507, 
    81.59199, 82.02757, 82.41193, 82.73427, 82.98342, 83.1489, 83.22219, 
    83.19816, 83.07582, 82.85847, 82.55286, 82.16798, 81.71375, 81.19992, 
    80.63553, 80.02852, 79.3857, 78.7128, 78.01461, 77.29511, 76.55762, 
    75.80494, 75.03938, 74.26292, 73.47726, 72.68385, 71.88396, 71.07871, 
    70.26908, 69.45595, 68.64011, 67.8223, 67.00318, 66.18338, 65.36349, 
    64.54404, 63.7256, 62.90866, 62.09375, 61.28136, 60.472, 59.66619, 
    58.86449, 58.06747, 57.27575, 56.49005, 55.71118, 54.94013, 54.17815, 
    53.42694, 52.68894, 51.96816, 51.27207, 50.61779, 50.05792, 49.78856,
  50.13831, 49.82203, 50.13831, 50.73761, 51.41262, 52.12174, 52.85207, 
    53.59786, 54.35592, 55.12421, 55.90129, 56.68607, 57.47766, 58.27533, 
    59.07841, 59.88634, 60.69857, 61.51461, 62.33397, 63.15618, 63.98077, 
    64.80728, 65.63524, 66.46416, 67.29355, 68.12287, 68.95158, 69.77908, 
    70.60473, 71.42783, 72.2476, 73.06319, 73.87363, 74.67781, 75.47445, 
    76.26205, 77.03884, 77.80273, 78.55116, 79.28102, 79.9885, 80.66886, 
    81.31624, 81.92336, 82.48131, 82.97943, 83.40544, 83.7461, 83.98865, 
    84.12289, 84.14357, 84.05181, 83.85507, 83.56548, 83.19739, 82.76532, 
    82.28255, 81.76051, 81.20869, 80.63488, 80.04536, 79.44525, 78.83873, 
    78.22928, 77.61981, 77.01285, 76.41058, 75.81495, 75.22776, 74.65067, 
    74.08529, 73.53316, 72.99581, 72.47482, 71.97176, 71.48833, 71.02627, 
    70.58746, 70.17387, 69.78767, 69.43108, 69.10648, 68.81618, 68.56233, 
    68.34651, 68.16934, 68.0299, 67.92546, 67.85175, 67.80377, 67.77703, 
    67.76848, 67.77703, 67.80377, 67.85175, 67.92546, 68.0299, 68.16934, 
    68.34651, 68.56233, 68.81618, 69.10648, 69.43108, 69.78767, 70.17387, 
    70.58746, 71.02627, 71.48833, 71.97176, 72.47482, 72.99581, 73.53316, 
    74.08529, 74.65067, 75.22776, 75.81495, 76.41058, 77.01285, 77.61981, 
    78.22928, 78.83873, 79.44525, 80.04536, 80.63488, 81.20869, 81.76051, 
    82.28255, 82.76532, 83.19739, 83.56548, 83.85507, 84.05181, 84.14357, 
    84.12289, 83.98865, 83.7461, 83.40544, 82.97943, 82.48131, 81.92336, 
    81.31624, 80.66886, 79.9885, 79.28102, 78.55116, 77.80273, 77.03884, 
    76.26205, 75.47445, 74.67781, 73.87363, 73.06319, 72.2476, 71.42783, 
    70.60473, 69.77908, 68.95158, 68.12287, 67.29355, 66.46416, 65.63524, 
    64.80728, 63.98077, 63.15618, 62.33397, 61.51461, 60.69857, 59.88634, 
    59.07841, 58.27533, 57.47766, 56.68607, 55.90129, 55.12421, 54.35592, 
    53.59786, 52.85207, 52.12174, 51.41262, 50.73761, 50.13831, 49.82203,
  50.22058, 49.85293, 50.22058, 50.85079, 51.54044, 52.2587, 52.99587, 
    53.7474, 54.51064, 55.28381, 56.06565, 56.85516, 57.65152, 58.45404, 
    59.26212, 60.07522, 60.89283, 61.71447, 62.5397, 63.36809, 64.19919, 
    65.03258, 65.86784, 66.70451, 67.54215, 68.3803, 69.21847, 70.05612, 
    70.89272, 71.72765, 72.56026, 73.3898, 74.21546, 75.0363, 75.85124, 
    76.65901, 77.45811, 78.24673, 79.02264, 79.7831, 80.52465, 81.24287, 
    81.93207, 82.58489, 83.19183, 83.7407, 84.21644, 84.60144, 84.8773, 
    85.02817, 85.0452, 84.92979, 84.69338, 84.35401, 83.93176, 83.44546, 
    82.91103, 82.34128, 81.74622, 81.13358, 80.50941, 79.87843, 79.24444, 
    78.61051, 77.97923, 77.35279, 76.73311, 76.12192, 75.52081, 74.93131, 
    74.35487, 73.79295, 73.24699, 72.71852, 72.20911, 71.72043, 71.25428, 
    70.8126, 70.39751, 70.01136, 69.65664, 69.33606, 69.05238, 68.80817, 
    68.60532, 68.44429, 68.32323, 68.23756, 68.18073, 68.14582, 68.1272, 
    68.12138, 68.1272, 68.14582, 68.18073, 68.23756, 68.32323, 68.44429, 
    68.60532, 68.80817, 69.05238, 69.33606, 69.65664, 70.01136, 70.39751, 
    70.8126, 71.25428, 71.72043, 72.20911, 72.71852, 73.24699, 73.79295, 
    74.35487, 74.93131, 75.52081, 76.12192, 76.73311, 77.35279, 77.97923, 
    78.61051, 79.24444, 79.87843, 80.50941, 81.13358, 81.74622, 82.34128, 
    82.91103, 83.44546, 83.93176, 84.35401, 84.69338, 84.92979, 85.0452, 
    85.02817, 84.8773, 84.60144, 84.21644, 83.7407, 83.19183, 82.58489, 
    81.93207, 81.24287, 80.52465, 79.7831, 79.02264, 78.24673, 77.45811, 
    76.65901, 75.85124, 75.0363, 74.21546, 73.3898, 72.56026, 71.72765, 
    70.89272, 70.05612, 69.21847, 68.3803, 67.54215, 66.70451, 65.86784, 
    65.03258, 64.19919, 63.36809, 62.5397, 61.71447, 60.89283, 60.07522, 
    59.26212, 58.45404, 57.65152, 56.85516, 56.06565, 55.28381, 54.51064, 
    53.7474, 52.99587, 52.2587, 51.54044, 50.85079, 50.22058, 49.85293,
  50.30153, 49.88158, 50.30153, 50.95307, 51.6522, 52.37652, 53.11841, 
    53.87404, 54.64109, 55.41796, 56.20347, 56.99667, 57.7968, 58.60321, 
    59.41531, 60.23259, 61.05458, 61.88081, 62.71086, 63.54433, 64.38081, 
    65.21989, 66.06121, 66.90434, 67.74889, 68.59444, 69.44056, 70.28679, 
    71.13266, 71.97765, 72.82121, 73.66272, 74.50151, 75.33682, 76.16777, 
    76.99332, 77.81229, 78.62318, 79.42419, 80.21306, 80.98686, 81.74178, 
    82.47274, 83.17283, 83.83259, 84.439, 84.97443, 85.41604, 85.73708, 
    85.91196, 85.92498, 85.77793, 85.48977, 85.08855, 84.60263, 84.05585, 
    83.46651, 82.84804, 82.21024, 81.5603, 80.90357, 80.24413, 79.5852, 
    78.92934, 78.2787, 77.63513, 77.00027, 76.37559, 75.7625, 75.16235, 
    74.57648, 74.00624, 73.45302, 72.91828, 72.40358, 71.91061, 71.44122, 
    70.99744, 70.58155, 70.19614, 69.84407, 69.52856, 69.25304, 69.02085, 
    68.83453, 68.69438, 68.59689, 68.53433, 68.4969, 68.47589, 68.46538, 
    68.4622, 68.46538, 68.47589, 68.4969, 68.53433, 68.59689, 68.69438, 
    68.83453, 69.02085, 69.25304, 69.52856, 69.84407, 70.19614, 70.58155, 
    70.99744, 71.44122, 71.91061, 72.40358, 72.91828, 73.45302, 74.00624, 
    74.57648, 75.16235, 75.7625, 76.37559, 77.00027, 77.63513, 78.2787, 
    78.92934, 79.5852, 80.24413, 80.90357, 81.5603, 82.21024, 82.84804, 
    83.46651, 84.05585, 84.60263, 85.08855, 85.48977, 85.77793, 85.92498, 
    85.91196, 85.73708, 85.41604, 84.97443, 84.439, 83.83259, 83.17283, 
    82.47274, 81.74178, 80.98686, 80.21306, 79.42419, 78.62318, 77.81229, 
    76.99332, 76.16777, 75.33682, 74.50151, 73.66272, 72.82121, 71.97765, 
    71.13266, 70.28679, 69.44056, 68.59444, 67.74889, 66.90434, 66.06121, 
    65.21989, 64.38081, 63.54433, 62.71086, 61.88081, 61.05458, 60.23259, 
    59.41531, 58.60321, 57.7968, 56.99667, 56.20347, 55.41796, 54.64109, 
    53.87404, 53.11841, 52.37652, 51.6522, 50.95307, 50.30153, 49.88158,
  50.37637, 49.90826, 50.37637, 51.04055, 51.74527, 52.47337, 53.21838, 
    53.97686, 54.74664, 55.52623, 56.31447, 57.11048, 57.91351, 58.72291, 
    59.53815, 60.3587, 61.18411, 62.01395, 62.84782, 63.68532, 64.52607, 
    65.36971, 66.21586, 67.06417, 67.91426, 68.76576, 69.61829, 70.47145, 
    71.32484, 72.17802, 73.03053, 73.88186, 74.73148, 75.57877, 76.42307, 
    77.26357, 78.09936, 78.92931, 79.75209, 80.56596, 81.36869, 82.15731, 
    82.92773, 83.67418, 84.38824, 85.0574, 85.6628, 86.17659, 86.56061, 
    86.77191, 86.78035, 86.58852, 86.23083, 85.75279, 85.19376, 84.58217, 
    83.93718, 83.2715, 82.59374, 81.90987, 81.22417, 80.53986, 79.85943, 
    79.18487, 78.5179, 77.85999, 77.21249, 76.57664, 75.95368, 75.3448, 
    74.75121, 74.17419, 73.61507, 73.07526, 72.55632, 72.05994, 71.58805, 
    71.14278, 70.72661, 70.34241, 69.99353, 69.68393, 69.41816, 69.20107, 
    69.0366, 68.92483, 68.85826, 68.82292, 68.80523, 68.79654, 68.79253, 
    68.79137, 68.79253, 68.79654, 68.80523, 68.82292, 68.85826, 68.92483, 
    69.0366, 69.20107, 69.41816, 69.68393, 69.99353, 70.34241, 70.72661, 
    71.14278, 71.58805, 72.05994, 72.55632, 73.07526, 73.61507, 74.17419, 
    74.75121, 75.3448, 75.95368, 76.57664, 77.21249, 77.85999, 78.5179, 
    79.18487, 79.85943, 80.53986, 81.22417, 81.90987, 82.59374, 83.2715, 
    83.93718, 84.58217, 85.19376, 85.75279, 86.23083, 86.58852, 86.78035, 
    86.77191, 86.56061, 86.17659, 85.6628, 85.0574, 84.38824, 83.67418, 
    82.92773, 82.15731, 81.36869, 80.56596, 79.75209, 78.92931, 78.09936, 
    77.26357, 76.42307, 75.57877, 74.73148, 73.88186, 73.03053, 72.17802, 
    71.32484, 70.47145, 69.61829, 68.76576, 67.91426, 67.06417, 66.21586, 
    65.36971, 64.52607, 63.68532, 62.84782, 62.01395, 61.18411, 60.3587, 
    59.53815, 58.72291, 57.91351, 57.11048, 56.31447, 55.52623, 54.74664, 
    53.97686, 53.21838, 52.47337, 51.74527, 51.04055, 50.37637, 49.90826,
  50.43979, 49.93322, 50.43979, 51.11018, 51.81787, 52.54819, 53.29517, 
    54.05554, 54.82721, 55.6087, 56.39891, 57.19695, 58.00209, 58.8137, 
    59.63124, 60.45423, 61.2822, 62.11474, 62.95146, 63.79198, 64.63595, 
    65.48301, 66.33281, 67.18504, 68.03931, 68.89533, 69.75274, 70.61118, 
    71.47032, 72.32977, 73.18914, 74.04804, 74.90604, 75.76264, 76.61736, 
    77.4696, 78.3187, 79.16389, 80.00422, 80.83852, 81.66531, 82.48254, 
    83.28741, 84.07583, 84.8415, 85.57432, 86.25728, 86.86075, 87.33431, 
    87.60472, 87.60763, 87.34742, 86.89431, 86.3233, 85.68491, 85.00868, 
    84.31155, 83.60366, 82.89138, 82.17895, 81.46935, 80.76483, 80.06713, 
    79.37772, 78.69786, 78.02872, 77.37135, 76.72684, 76.09622, 75.48059, 
    74.88106, 74.29882, 73.73515, 73.19144, 72.66924, 72.17028, 71.6965, 
    71.2502, 70.83404, 70.45123, 70.10575, 69.80266, 69.54853, 69.35167, 
    69.22012, 69.15179, 69.12489, 69.11536, 69.11171, 69.11018, 69.10952, 
    69.10934, 69.10952, 69.11018, 69.11171, 69.11536, 69.12489, 69.15179, 
    69.22012, 69.35167, 69.54853, 69.80266, 70.10575, 70.45123, 70.83404, 
    71.2502, 71.6965, 72.17028, 72.66924, 73.19144, 73.73515, 74.29882, 
    74.88106, 75.48059, 76.09622, 76.72684, 77.37135, 78.02872, 78.69786, 
    79.37772, 80.06713, 80.76483, 81.46935, 82.17895, 82.89138, 83.60366, 
    84.31155, 85.00868, 85.68491, 86.3233, 86.89431, 87.34742, 87.60763, 
    87.60472, 87.33431, 86.86075, 86.25728, 85.57432, 84.8415, 84.07583, 
    83.28741, 82.48254, 81.66531, 80.83852, 80.00422, 79.16389, 78.3187, 
    77.4696, 76.61736, 75.76264, 74.90604, 74.04804, 73.18914, 72.32977, 
    71.47032, 70.61118, 69.75274, 68.89533, 68.03931, 67.18504, 66.33281, 
    65.48301, 64.63595, 63.79198, 62.95146, 62.11474, 61.2822, 60.45423, 
    59.63124, 58.8137, 58.00209, 57.19695, 56.39891, 55.6087, 54.82721, 
    54.05554, 53.29517, 52.54819, 51.81787, 51.11018, 50.43979, 49.93322,
  50.48727, 49.9567, 50.48727, 51.16006, 51.86916, 52.60069, 53.34884, 
    54.11039, 54.88327, 55.666, 56.45752, 57.25692, 58.06347, 58.87658, 
    59.6957, 60.52034, 61.35005, 62.18444, 63.02311, 63.8657, 64.71188, 
    65.56129, 66.41361, 67.26852, 68.1257, 68.98485, 69.84563, 70.70774, 
    71.57086, 72.43467, 73.29884, 74.16303, 75.02689, 75.89005, 76.75213, 
    77.61269, 78.47128, 79.3274, 80.18045, 81.02972, 81.87433, 82.71316, 
    83.54466, 84.36656, 85.17532, 85.96491, 86.72411, 87.42961, 88.02856, 
    88.40409, 88.39936, 88.02417, 87.44224, 86.76824, 86.05346, 85.32051, 
    84.58044, 83.83923, 83.10052, 82.3667, 81.63949, 80.92026, 80.21013, 
    79.51008, 78.82105, 78.14394, 77.47961, 76.82898, 76.19297, 75.57259, 
    74.96886, 74.38295, 73.81608, 73.2696, 72.74509, 72.24426, 71.76914, 
    71.32211, 70.906, 70.52443, 70.1821, 69.88578, 69.64649, 69.48528, 
    69.42566, 69.41785, 69.41682, 69.4166, 69.41654, 69.41651, 69.4165, 
    69.4165, 69.4165, 69.41651, 69.41654, 69.4166, 69.41682, 69.41785, 
    69.42566, 69.48528, 69.64649, 69.88578, 70.1821, 70.52443, 70.906, 
    71.32211, 71.76914, 72.24426, 72.74509, 73.2696, 73.81608, 74.38295, 
    74.96886, 75.57259, 76.19297, 76.82898, 77.47961, 78.14394, 78.82105, 
    79.51008, 80.21013, 80.92026, 81.63949, 82.3667, 83.10052, 83.83923, 
    84.58044, 85.32051, 86.05346, 86.76824, 87.44224, 88.02417, 88.39936, 
    88.40409, 88.02856, 87.42961, 86.72411, 85.96491, 85.17532, 84.36656, 
    83.54466, 82.71316, 81.87433, 81.02972, 80.18045, 79.3274, 78.47128, 
    77.61269, 76.75213, 75.89005, 75.02689, 74.16303, 73.29884, 72.43467, 
    71.57086, 70.70774, 69.84563, 68.98485, 68.1257, 67.26852, 66.41361, 
    65.56129, 64.71188, 63.8657, 63.02311, 62.18444, 61.35005, 60.52034, 
    59.6957, 58.87658, 58.06347, 57.25692, 56.45752, 55.666, 54.88327, 
    54.11039, 53.34884, 52.60069, 51.86916, 51.16006, 50.48727, 49.9567,
  50.51608, 49.97889, 50.51608, 51.18951, 51.89921, 52.63133, 53.38007, 
    54.14225, 54.91582, 55.69927, 56.49147, 57.29165, 58.09902, 58.91298, 
    59.73299, 60.55857, 61.38928, 62.22474, 63.06453, 63.90832, 64.75574, 
    65.6065, 66.46028, 67.31674, 68.17557, 69.03654, 69.89927, 70.76348, 
    71.62891, 72.49525, 73.36219, 74.22945, 75.09672, 75.96371, 76.83007, 
    77.69551, 78.55972, 79.42227, 80.28288, 81.14109, 81.99649, 82.84852, 
    83.69659, 84.5398, 85.37699, 86.20615, 87.02346, 87.82003, 88.56853, 
    89.14749, 89.12862, 88.54444, 87.81496, 87.05143, 86.27943, 85.50751, 
    84.73938, 83.97713, 83.22209, 82.47529, 81.7375, 81.00948, 80.29199, 
    79.58566, 78.89123, 78.20946, 77.54105, 76.88683, 76.24767, 75.6245, 
    75.01831, 74.43027, 73.86143, 73.3133, 72.78741, 72.28542, 71.80939, 
    71.36184, 70.94566, 70.56478, 70.22474, 69.93495, 69.72819, 69.71326, 
    69.71326, 69.71326, 69.71326, 69.71326, 69.71326, 69.71326, 69.71326, 
    69.71326, 69.71326, 69.71326, 69.71326, 69.71326, 69.71326, 69.71326, 
    69.71326, 69.71326, 69.72819, 69.93495, 70.22474, 70.56478, 70.94566, 
    71.36184, 71.80939, 72.28542, 72.78741, 73.3133, 73.86143, 74.43027, 
    75.01831, 75.6245, 76.24767, 76.88683, 77.54105, 78.20946, 78.89123, 
    79.58566, 80.29199, 81.00948, 81.7375, 82.47529, 83.22209, 83.97713, 
    84.73938, 85.50751, 86.27943, 87.05143, 87.81496, 88.54444, 89.12862, 
    89.14749, 88.56853, 87.82003, 87.02346, 86.20615, 85.37699, 84.5398, 
    83.69659, 82.84852, 81.99649, 81.14109, 80.28288, 79.42227, 78.55972, 
    77.69551, 76.83007, 75.96371, 75.09672, 74.22945, 73.36219, 72.49525, 
    71.62891, 70.76348, 69.89927, 69.03654, 68.17557, 67.31674, 66.46028, 
    65.6065, 64.75574, 63.90832, 63.06453, 62.22474, 61.38928, 60.55857, 
    59.73299, 58.91298, 58.09902, 57.29165, 56.49147, 55.69927, 54.91582, 
    54.14225, 53.38007, 52.63133, 51.89921, 51.18951, 50.51608, 49.97889,
  50.52546, 50, 50.52546, 51.19905, 51.90889, 52.64119, 53.39014, 54.15252, 
    54.92627, 55.70993, 56.5024, 57.30281, 58.11044, 58.92467, 59.74496, 
    60.57084, 61.40187, 62.23765, 63.0778, 63.92197, 64.76981, 65.62101, 
    66.47523, 67.33219, 68.19157, 69.05309, 69.91644, 70.78135, 71.64751, 
    72.51466, 73.38249, 74.25074, 75.1191, 75.9873, 76.85506, 77.72208, 
    78.58806, 79.45272, 80.31577, 81.17689, 82.03579, 82.89217, 83.74571, 
    84.5961, 85.44302, 86.28614, 87.12513, 87.95965, 88.78936, 89.6139, 
    89.56709, 88.75397, 87.94714, 87.14697, 86.35389, 85.5683, 84.79064, 
    84.02137, 83.26095, 82.50986, 81.76862, 81.03777, 80.31787, 79.60953, 
    78.91336, 78.23006, 77.56034, 76.90497, 76.26479, 75.64072, 75.03372, 
    74.44492, 73.87549, 73.3268, 72.80037, 72.29797, 71.82161, 71.37377, 
    70.95746, 70.57668, 70.23724, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 
    70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70.23724, 70.57668, 70.95746, 
    71.37377, 71.82161, 72.29797, 72.80037, 73.3268, 73.87549, 74.44492, 
    75.03372, 75.64072, 76.26479, 76.90497, 77.56034, 78.23006, 78.91336, 
    79.60953, 80.31787, 81.03777, 81.76862, 82.50986, 83.26095, 84.02137, 
    84.79064, 85.5683, 86.35389, 87.14697, 87.94714, 88.75397, 89.56709, 
    89.6139, 88.78936, 87.95965, 87.12513, 86.28614, 85.44302, 84.5961, 
    83.74571, 82.89217, 82.03579, 81.17689, 80.31577, 79.45272, 78.58806, 
    77.72208, 76.85506, 75.9873, 75.1191, 74.25074, 73.38249, 72.51466, 
    71.64751, 70.78135, 69.91644, 69.05309, 68.19157, 67.33219, 66.47523, 
    65.62101, 64.76981, 63.92197, 63.0778, 62.23765, 61.40187, 60.57084, 
    59.74496, 58.92467, 58.11044, 57.30281, 56.5024, 55.70993, 54.92627, 
    54.15252, 53.39014, 52.64119, 51.90889, 51.19905, 50.52546, 50,
  50.51608, 49.97889, 50.51608, 51.18951, 51.89921, 52.63133, 53.38007, 
    54.14225, 54.91582, 55.69927, 56.49147, 57.29165, 58.09902, 58.91298, 
    59.73299, 60.55857, 61.38928, 62.22474, 63.06453, 63.90832, 64.75574, 
    65.6065, 66.46028, 67.31674, 68.17557, 69.03654, 69.89927, 70.76348, 
    71.62891, 72.49525, 73.36219, 74.22945, 75.09672, 75.96371, 76.83007, 
    77.69551, 78.55972, 79.42227, 80.28288, 81.14109, 81.99649, 82.84852, 
    83.69659, 84.5398, 85.37699, 86.20615, 87.02346, 87.82003, 88.56853, 
    89.14749, 89.12862, 88.54444, 87.81496, 87.05143, 86.27943, 85.50751, 
    84.73938, 83.97713, 83.22209, 82.47529, 81.7375, 81.00948, 80.29199, 
    79.58566, 78.89123, 78.20946, 77.54105, 76.88683, 76.24767, 75.6245, 
    75.01831, 74.43027, 73.86143, 73.3133, 72.78741, 72.28542, 71.80939, 
    71.36184, 70.94566, 70.56478, 70.22474, 69.93495, 69.72819, 69.71326, 
    69.71326, 69.71326, 69.71326, 69.71326, 69.71326, 69.71326, 69.71326, 
    69.71326, 69.71326, 69.71326, 69.71326, 69.71326, 69.71326, 69.71326, 
    69.71326, 69.71326, 69.72819, 69.93495, 70.22474, 70.56478, 70.94566, 
    71.36184, 71.80939, 72.28542, 72.78741, 73.3133, 73.86143, 74.43027, 
    75.01831, 75.6245, 76.24767, 76.88683, 77.54105, 78.20946, 78.89123, 
    79.58566, 80.29199, 81.00948, 81.7375, 82.47529, 83.22209, 83.97713, 
    84.73938, 85.50751, 86.27943, 87.05143, 87.81496, 88.54444, 89.12862, 
    89.14749, 88.56853, 87.82003, 87.02346, 86.20615, 85.37699, 84.5398, 
    83.69659, 82.84852, 81.99649, 81.14109, 80.28288, 79.42227, 78.55972, 
    77.69551, 76.83007, 75.96371, 75.09672, 74.22945, 73.36219, 72.49525, 
    71.62891, 70.76348, 69.89927, 69.03654, 68.17557, 67.31674, 66.46028, 
    65.6065, 64.75574, 63.90832, 63.06453, 62.22474, 61.38928, 60.55857, 
    59.73299, 58.91298, 58.09902, 57.29165, 56.49147, 55.69927, 54.91582, 
    54.14225, 53.38007, 52.63133, 51.89921, 51.18951, 50.51608, 49.97889 ;

 nav_lon =
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, -3.999688, -1.999661, 0.0003655546, 2.000391, 4.000415, 
    6.000439, 8.000461, 10.00048, 12.0005, 14.00052, 16.00053, 18.00055, 
    20.00056, 22.00057, 24.00057, 26.00058, 28.00058, 30.00058, 32.00058, 
    34.00058, 36.00057, 38.00056, 40.00055, 42.00054, 44.00053, 46.00051, 
    48.00049, 50.00047, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 
    62.00031, 64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 
    76.00008, 78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, 26.50045, 27.50045, 28.50045, 29.50045, 30.50045, 31.50045, 
    32.50045, 33.50045, 34.50045, 35.50045, 36.48142, 37.4082, 38.25387, 
    39.00387, 39.6582, 40.23142, 40.75045, 41.25045, 41.75045, 42.25045, 
    42.75045, 43.25045, 43.80754, 44.52721, 45.4902, 46.7402, 48.27721, 
    50.05754, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 62.00031, 
    64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 76.00008, 
    78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, 26.50045, 27.50045, 28.50045, 29.50045, 30.50045, 31.50045, 
    32.50045, 33.50045, 34.50045, 35.50045, 36.48142, 37.4082, 38.25387, 
    39.00387, 39.6582, 40.23142, 40.75045, 41.25045, 41.75045, 42.25045, 
    42.75045, 43.25045, 43.80754, 44.52721, 45.4902, 46.7402, 48.27721, 
    50.05754, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 62.00031, 
    64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 76.00008, 
    78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, 26.50045, 27.50045, 28.50045, 29.50045, 30.50045, 31.50045, 
    32.50045, 33.50045, 34.50045, 35.50045, 36.48142, 37.4082, 38.25387, 
    39.00387, 39.6582, 40.23142, 40.75045, 41.25045, 41.75045, 42.25045, 
    42.75045, 43.25045, 43.80754, 44.52721, 45.4902, 46.7402, 48.27721, 
    50.05754, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 62.00031, 
    64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 76.00008, 
    78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, 26.50045, 27.50045, 28.50045, 29.50045, 30.50045, 31.50045, 
    32.50045, 33.50045, 34.50045, 35.50045, 36.48142, 37.4082, 38.25387, 
    39.00387, 39.6582, 40.23142, 40.75045, 41.25045, 41.75045, 42.25045, 
    42.75045, 43.25045, 43.80754, 44.52721, 45.4902, 46.7402, 48.27721, 
    50.05754, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 62.00031, 
    64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 76.00008, 
    78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, 26.50045, 27.50045, 28.50045, 29.50045, 30.50045, 31.50045, 
    32.50045, 33.50045, 34.50045, 35.50045, 36.48142, 37.4082, 38.25387, 
    39.00387, 39.6582, 40.23142, 40.75045, 41.25045, 41.75045, 42.25045, 
    42.75045, 43.25045, 43.80754, 44.52721, 45.4902, 46.7402, 48.27721, 
    50.05754, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 62.00031, 
    64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 76.00008, 
    78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, 26.50045, 27.50045, 28.50045, 29.50045, 30.50045, 31.50045, 
    32.50045, 33.50045, 34.50045, 35.50045, 36.48142, 37.4082, 38.25387, 
    39.00387, 39.6582, 40.23142, 40.75045, 41.25045, 41.75045, 42.25045, 
    42.75045, 43.25045, 43.80754, 44.52721, 45.4902, 46.7402, 48.27721, 
    50.05754, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 62.00031, 
    64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 76.00008, 
    78.00004, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, 26.50045, 27.50045, 28.50045, 29.50045, 30.50045, 31.50045, 
    32.50045, 33.50045, 34.50045, 35.50045, 36.48142, 37.4082, 38.25387, 
    39.00387, 39.6582, 40.23142, 40.75045, 41.25045, 41.75045, 42.25045, 
    42.75045, 43.25045, 43.80754, 44.52721, 45.4902, 46.7402, 48.27721, 
    50.05754, 52.00045, 54.00043, 56.0004, 58.00037, 60.00034, 62.00031, 
    64.00028, 66.00025, 68.00021, 70.00018, 72.00014, 74.00011, 76.00008, 
    78.00004, 80,
  78, 80, 82, 84, 86, 88, 90, 92, 94, 96, 98, 100, 102, 104, 106, 108, 110, 
    112, 114, 116, 118, 120, 122, 124, 126, 128, 130, 132, 134, 136, 138, 
    140, 142, 144, 146, 148, 150, 152, 154, 156, 158, 160, 162, 164, 166, 
    168, 170, 172, 174, 176, 178, 180, -178, -176, -174, -172, -170, -168, 
    -166, -164, -162, -160, -158, -156, -154, -152, -150, -148, -146, -144, 
    -142, -140, -138, -136, -134, -132, -130, -128, -126, -124, -122, -120, 
    -118, -116, -114, -112, -110, -108, -106, -104, -102, -100, -98, -96, 
    -94, -92, -90, -88, -86, -84, -82, -80, -78, -76, -74, -72, -70, -68, 
    -66, -64, -62, -60, -58, -56, -54, -52, -50, -48, -46, -44, -42, -40, 
    -38, -36, -34, -32, -30, -28, -26, -24, -22, -20, -18, -16, -14, -12, 
    -10, -8, -6, 26.5, 27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 
    36.48097, 37.40775, 38.25342, 39.00342, 39.65775, 40.23097, 40.75, 41.25, 
    41.75, 42.25, 42.75, 43.25, 43.80709, 44.52676, 45.48975, 46.73975, 
    48.27676, 50.05709, 52, 54, 56, 58, 60, 62, 64, 66, 68, 70, 72, 74, 76, 
    78, 80,
  78.00001, 80, 81.99999, 83.99999, 85.99998, 87.99998, 89.99998, 91.99998, 
    93.99997, 95.99997, 97.99996, 99.99996, 102, 104, 106, 107.9999, 
    109.9999, 111.9999, 113.9999, 115.9999, 117.9999, 119.9999, 121.9999, 
    123.9999, 125.9999, 127.9999, 129.9999, 131.9999, 133.9999, 135.9999, 
    137.9999, 139.9999, 141.9999, 143.9999, 145.9999, 147.9999, 149.9999, 
    152, 154, 156, 158, 160, 162, 164, 166, 168, 170, 172, 174, 176, 178, 
    180, -178, -176, -174, -172, -170, -168, -166, -164, -162, -160, -158, 
    -156, -154, -152, -150, -148, -146, -144, -142, -140, -138, -136, -134, 
    -132, -130, -128, -126, -124, -122, -120, -118, -116, -114, -112, -110, 
    -108, -106, -104, -102, -100, -98, -96.00001, -94.00001, -92.00001, 
    -90.00002, -88.00002, -86.00002, -84.00002, -82.00002, -80.00002, 
    -78.00002, -76.00002, -74.00002, -72.00003, -70.00003, -68.00003, 
    -66.00003, -64.00003, -62.00003, -60.00003, -58.00003, -56.00003, 
    -54.00003, -52.00003, -50.00003, -48.00003, -46.00002, -44.00002, 
    -42.00002, -40.00002, -38.00002, -36.00002, -34.00001, -32.00001, 
    -30.00001, -28, -26, -24, -21.99999, -19.99999, -17.99999, -15.99998, 
    -13.99998, -11.99998, -9.999974, -7.999971, -5.999968, 26.50005, 
    27.50005, 28.50005, 29.50005, 30.50005, 31.50005, 32.50005, 33.50005, 
    34.50005, 35.50005, 36.48102, 37.4078, 38.25347, 39.00347, 39.6578, 
    40.23102, 40.75005, 41.25005, 41.75005, 42.25005, 42.75005, 43.25005, 
    43.80714, 44.52681, 45.4898, 46.7398, 48.27681, 50.05714, 52.00005, 
    54.00005, 56.00005, 58.00004, 60.00004, 62.00003, 64.00003, 66.00003, 
    68.00002, 70.00002, 72.00002, 74.00002, 76.00001, 78.00001, 80,
  78.00004, 80, 81.99996, 83.99992, 85.99989, 87.99986, 89.99982, 91.99979, 
    93.99975, 95.99972, 97.99969, 99.99966, 101.9996, 103.9996, 105.9996, 
    107.9995, 109.9995, 111.9995, 113.9995, 115.9995, 117.9995, 119.9994, 
    121.9994, 123.9994, 125.9994, 127.9994, 129.9994, 131.9994, 133.9994, 
    135.9994, 137.9994, 139.9995, 141.9995, 143.9995, 145.9995, 147.9995, 
    149.9995, 151.9995, 153.9996, 155.9996, 157.9996, 159.9996, 161.9997, 
    163.9997, 165.9997, 167.9997, 169.9998, 171.9998, 173.9998, 175.9999, 
    177.9999, 179.9999, -178, -176, -174, -172, -169.9999, -167.9999, 
    -165.9999, -163.9999, -161.9998, -159.9998, -157.9998, -155.9998, 
    -153.9998, -151.9998, -149.9998, -147.9998, -145.9997, -143.9997, 
    -141.9997, -139.9997, -137.9997, -135.9997, -133.9997, -131.9997, 
    -129.9998, -127.9998, -125.9998, -123.9998, -121.9998, -119.9998, 
    -117.9998, -115.9998, -113.9999, -111.9999, -109.9999, -107.9999, 
    -105.9999, -104, -102, -100, -98.00002, -96.00005, -94.00006, -92.00008, 
    -90.00011, -88.00012, -86.00014, -84.00016, -82.00018, -80.00019, 
    -78.00021, -76.00022, -74.00023, -72.00024, -70.00025, -68.00026, 
    -66.00026, -64.00027, -62.00027, -60.00027, -58.00027, -56.00026, 
    -54.00026, -52.00025, -50.00024, -48.00023, -46.00022, -44.0002, 
    -42.00019, -40.00017, -38.00015, -36.00013, -34.00011, -32.00008, 
    -30.00006, -28.00003, -26.00001, -23.99998, -21.99995, -19.99992, 
    -17.99989, -15.99986, -13.99983, -11.9998, -9.999774, -7.999745, 
    -5.999716, 26.50045, 27.50045, 28.50045, 29.50045, 30.50045, 31.50045, 
    32.50045, 33.50045, 34.50045, 35.50045, 36.48142, 37.4082, 38.25387, 
    39.00387, 8.530076, 9.530076, 10.53008, 11.53008, 12.53008, 13.53008, 
    14.53008, 15.53008, 16.53008, 17.53008, 18.53008, 19.53008, 20.53008, 
    21.53008, 22.53008, 23.53008, 24.53008, 58.00004, 60.00004, 62.00003, 
    64.00003, 66.00003, 68.00002, 70.00002, 32.53008, 33.53008, 34.53008, 
    35.53008, 80,
  78.00014, 80, 81.99986, 83.99971, 85.99957, 87.99944, 89.9993, 91.99916, 
    93.99903, 95.9989, 97.99878, 99.99866, 101.9985, 103.9984, 105.9983, 
    107.9982, 109.9982, 111.9981, 113.998, 115.9979, 117.9979, 119.9978, 
    121.9978, 123.9978, 125.9977, 127.9977, 129.9977, 131.9977, 133.9977, 
    135.9977, 137.9978, 139.9978, 141.9978, 143.9979, 145.998, 147.998, 
    149.9981, 151.9982, 153.9983, 155.9984, 157.9985, 159.9986, 161.9987, 
    163.9988, 165.9989, 167.999, 169.9991, 171.9992, 173.9993, 175.9995, 
    177.9996, 179.9997, -178.0002, -176.0001, -174, -171.9999, -169.9998, 
    -167.9997, -165.9996, -163.9995, -161.9994, -159.9993, -157.9993, 
    -155.9992, -153.9991, -151.9991, -149.9991, -147.999, -145.999, -143.999, 
    -141.9989, -139.9989, -137.9989, -135.9989, -133.999, -131.999, -129.999, 
    -127.999, -125.9991, -123.9991, -121.9992, -119.9992, -117.9993, 
    -115.9994, -113.9994, -111.9995, -109.9996, -107.9997, -105.9997, 
    -103.9998, -101.9999, -100, -98.00008, -96.00017, -94.00025, -92.00033, 
    -90.00041, -88.00049, -86.00056, -84.00063, -82.00069, -80.00076, 
    -78.00082, -76.00087, -74.00092, -72.00095, -70.00098, -68.00101, 
    -66.00104, -64.00105, -62.00106, -60.00106, -58.00105, -56.00104, 
    -54.00101, -52.00099, -50.00095, -48.00091, -46.00086, -44.0008, 
    -42.00074, -40.00066, -38.00059, -36.00051, -34.00042, -32.00033, 
    -30.00023, -28.00013, -26.00002, -23.99991, -21.9998, -19.99969, 
    -17.99957, -15.99946, -13.99934, -11.99923, -9.999109, -7.998994, 
    -5.998881, 26.50176, 27.50176, 28.50176, 29.50176, 30.50176, 31.50176, 
    32.50176, 33.50176, 34.50176, 35.50176, 36.48273, 37.4095, 38.25518, 
    39.00518, 8.530076, 9.530076, 10.53008, 11.53008, 12.53008, 13.53008, 
    14.53008, 15.53008, 16.53008, 17.53008, 18.53008, 19.53008, 20.53008, 
    21.53008, 22.53008, 23.53008, 24.53008, 25.53008, 26.53008, 27.53008, 
    28.53008, 29.53008, 30.53008, 31.53008, 32.53008, 33.53008, 34.53008, 
    35.53008, 80,
  78.00039, 80, 81.99961, 83.99922, 85.99884, 87.99846, 89.99809, 91.99772, 
    93.99737, 95.99702, 97.99668, 99.99636, 101.996, 103.9958, 105.9955, 
    107.9952, 109.995, 111.9948, 113.9946, 115.9944, 117.9942, 119.9941, 
    121.994, 123.9939, 125.9938, 127.9938, 129.9938, 131.9938, 133.9938, 
    135.9938, 137.9939, 139.994, 141.9941, 143.9943, 145.9944, 147.9946, 
    149.9948, 151.995, 153.9953, 155.9955, 157.9958, 159.996, 161.9963, 
    163.9966, 165.9969, 167.9972, 169.9976, 171.9979, 173.9982, 175.9985, 
    177.9988, 179.9991, -178.0005, -176.0002, -173.9999, -171.9996, 
    -169.9994, -167.9991, -165.9988, -163.9986, -161.9984, -159.9982, 
    -157.998, -155.9978, -153.9976, -151.9975, -149.9974, -147.9973, 
    -145.9972, -143.9971, -141.9971, -139.9971, -137.9971, -135.9971, 
    -133.9971, -131.9972, -129.9973, -127.9974, -125.9975, -123.9976, 
    -121.9978, -119.9979, -117.9981, -115.9983, -113.9985, -111.9987, 
    -109.9989, -107.9991, -105.9993, -103.9995, -101.9998, -100, -98.00023, 
    -96.00046, -94.00069, -92.00091, -90.00112, -88.00134, -86.00153, 
    -84.00172, -82.00191, -80.00208, -78.00224, -76.00237, -74.0025, 
    -72.00262, -70.00271, -68.00278, -66.00285, -64.00288, -62.00291, 
    -60.00291, -58.00289, -56.00285, -54.00279, -52.00271, -50.00262, 
    -48.00249, -46.00236, -44.0022, -42.00203, -40.00183, -38.00163, 
    -36.0014, -34.00116, -32.0009, -30.00064, -28.00036, -26.00007, 
    -23.99977, -21.99946, -19.99915, -17.99883, -15.99852, -13.99819, 
    -11.99787, -9.997556, -7.997241, -5.996931, 26.50478, 27.50478, 28.50478, 
    29.50478, 30.50478, 31.50478, 32.50478, 33.50176, 34.50176, 35.50176, 
    4.530076, 5.530076, 6.530076, 7.530076, 8.530076, 9.530076, 10.53008, 
    11.53008, 12.53008, 13.53008, 14.53008, 15.53008, 16.53008, 17.53008, 
    18.53008, 19.53008, 20.53008, 21.53008, 22.53008, 23.53008, 24.53008, 
    25.53008, 26.53008, 27.53008, 28.53008, 29.53008, 30.53008, 31.53008, 
    32.53008, 33.53008, 34.53008, 35.53008, 80,
  78.00085, 80, 81.99915, 83.99831, 85.99747, 87.99664, 89.99581, 91.99501, 
    93.99423, 95.99347, 97.99273, 99.99202, 101.9913, 103.9907, 105.9901, 
    107.9895, 109.989, 111.9885, 113.988, 115.9876, 117.9873, 119.987, 
    121.9867, 123.9865, 125.9864, 127.9863, 129.9862, 131.9862, 133.9863, 
    135.9864, 137.9865, 139.9867, 141.987, 143.9873, 145.9877, 147.9881, 
    149.9885, 151.989, 153.9895, 155.99, 157.9906, 159.9912, 161.9919, 
    163.9925, 165.9932, 167.9939, 169.9946, 171.9953, 173.996, 175.9967, 
    177.9974, 179.9981, -178.0012, -176.0005, -173.9998, -171.9992, 
    -169.9986, -167.998, -165.9974, -163.9969, -161.9964, -159.9959, 
    -157.9955, -155.9951, -153.9947, -151.9944, -149.9942, -147.9939, 
    -145.9938, -143.9936, -141.9936, -139.9935, -137.9935, -135.9936, 
    -133.9937, -131.9938, -129.994, -127.9942, -125.9944, -123.9947, 
    -121.995, -119.9954, -117.9958, -115.9962, -113.9966, -111.997, 
    -109.9975, -107.998, -105.9985, -103.999, -101.9995, -100, -98.00051, 
    -96.00102, -94.00153, -92.00201, -90.00249, -88.00296, -86.00341, 
    -84.00384, -82.00424, -80.00462, -78.00497, -76.00529, -74.00557, 
    -72.00582, -70.00603, -68.0062, -66.00634, -64.00642, -62.00648, 
    -60.00648, -58.00644, -56.00636, -54.00623, -52.00605, -50.00584, 
    -48.00557, -46.00526, -44.00492, -42.00453, -40.0041, -38.00363, 
    -36.00313, -34.00259, -32.00203, -30.00143, -28.00081, -26.00016, 
    -23.9995, -21.99881, -19.99812, -17.99741, -15.9967, -13.99599, 
    -11.99527, -9.994565, -7.993864, -5.993175, -3.992495, -4.469924, 
    -3.469924, -2.469924, -1.469924, -0.4699244, 0.5300756, 1.530076, 
    2.530076, 3.530076, 4.530076, 5.530076, 6.530076, 7.530076, 8.530076, 
    9.530076, 10.53008, 11.53008, 12.53008, 13.53008, 14.53008, 15.53008, 
    16.53008, 17.53008, 18.53008, 19.53008, 20.53008, 21.53008, 22.53008, 
    23.53008, 24.53008, 25.53008, 26.53008, 27.53008, 28.53008, 29.53008, 
    30.53008, 31.53008, 32.53008, 33.53008, 34.53008, 35.53008, 80,
  78.00162, 79.00162, 81.99838, 83.99678, 85.99518, 87.9936, 89.99204, 
    91.99052, 93.98902, 95.98757, 97.98616, 99.98481, 101.9835, 103.9823, 
    105.9811, 107.98, 109.979, 111.978, 113.9771, 115.9764, 117.9757, 
    119.9751, 121.9746, 123.9742, 125.9738, 127.9736, 129.9735, 131.9735, 
    133.9736, 135.9738, 137.9741, 139.9745, 141.9749, 143.9755, 145.9762, 
    147.9769, 149.9778, 151.9787, 153.9797, 155.9807, 157.9818, 159.983, 
    161.9842, 163.9855, 165.9868, 167.9881, 169.9895, 171.9909, 173.9922, 
    175.9936, 177.995, 179.9964, -178.0023, -176.0009, -173.9997, -171.9984, 
    -169.9972, -167.996, -165.9949, -163.9939, -161.9929, -159.992, 
    -157.9912, -155.9904, -153.9898, -151.9892, -149.9887, -147.9882, 
    -145.9879, -143.9877, -141.9875, -139.9874, -137.9874, -135.9875, 
    -133.9877, -131.988, -129.9883, -127.9887, -125.9892, -123.9898, 
    -121.9904, -119.9911, -117.9918, -115.9926, -113.9934, -111.9943, 
    -109.9952, -107.9961, -105.9971, -103.998, -101.999, -100, -98.00099, 
    -96.00197, -94.00294, -92.0039, -90.00483, -88.00573, -86.0066, 
    -84.00742, -82.0082, -80.00893, -78.00961, -76.01023, -74.01079, 
    -72.01127, -70.01168, -68.01202, -66.01228, -64.01247, -62.01256, 
    -60.01258, -58.0125, -56.01234, -54.0121, -52.01176, -50.01134, 
    -48.01083, -46.01024, -44.00957, -42.00882, -40.00798, -38.00708, 
    -36.0061, -34.00506, -32.00396, -30.0028, -28.00159, -26.00034, 
    -23.99905, -21.99772, -19.99637, -17.995, -15.99362, -13.99224, 
    -11.99085, -9.989478, -8.11004, -6.355933, -4.729666, -4.469924, 
    -3.469924, -2.469924, -1.469924, -0.4699244, 0.5300756, 1.530076, 
    2.530076, 3.530076, 4.530076, 5.530076, 6.530076, 7.530076, 8.530076, 
    9.530076, 10.53008, 11.53008, 12.53008, 13.53008, 14.53008, 15.53008, 
    16.53008, 17.53008, 18.53008, 19.53008, 20.53008, 21.53008, 22.53008, 
    23.53008, 24.53008, 25.53008, 26.53008, 27.53008, 28.53008, 29.53008, 
    30.53008, 31.53008, 32.53008, 33.53008, 34.53008, 35.53008, 36.53008,
  78.00277, 79.00162, 81.99723, 83.99446, 85.99172, 87.98901, 89.98633, 
    91.9837, 93.98112, 95.97862, 97.97619, 99.97384, 101.9716, 103.9694, 
    105.9674, 107.9655, 109.9637, 111.962, 113.9605, 115.9591, 117.9579, 
    119.9568, 121.9559, 123.9552, 125.9546, 127.9542, 129.9539, 131.9539, 
    133.954, 135.9543, 137.9548, 139.9554, 141.9563, 143.9572, 145.9584, 
    147.9597, 149.9611, 151.9627, 153.9644, 155.9662, 157.9681, 159.9702, 
    161.9723, 163.9745, 165.9768, 167.9792, 169.9815, 171.984, 173.9864, 
    175.9888, 177.9913, 179.9937, -178.004, -176.0016, -173.9994, -171.9971, 
    -169.995, -167.993, -165.991, -163.9892, -161.9875, -159.9859, -157.9844, 
    -155.9831, -153.9819, -151.9809, -149.98, -147.9793, -145.9787, 
    -143.9783, -141.978, -139.9779, -137.9779, -135.9781, -133.9784, 
    -131.9789, -129.9795, -127.9802, -125.9811, -123.982, -121.9831, 
    -119.9843, -117.9856, -115.987, -113.9884, -111.99, -109.9915, -107.9932, 
    -105.9948, -103.9965, -101.9983, -100, -98.00173, -96.00346, -94.00516, 
    -92.00683, -90.00846, -88.01004, -86.01156, -84.01302, -82.01439, 
    -80.01568, -78.01687, -76.01795, -74.01893, -72.01979, -70.02052, 
    -68.02113, -66.02159, -64.02191, -62.02209, -60.02213, -58.02201, 
    -56.02173, -54.02131, -52.02073, -50.01999, -48.0191, -46.01807, 
    -44.01689, -42.01556, -40.0141, -38.01251, -36.0108, -34.00896, 
    -32.00702, -30.00498, -28.00286, -26.00065, -23.99837, -21.99604, 
    -19.99366, -17.99125, -15.98882, -13.98639, -11.98396, -9.981542, -8.227, 
    -6.7231, -5.469924, -4.469924, -3.469924, -2.469924, -1.469924, 
    -0.4699244, 0.5300756, 1.530076, 2.530076, 3.530076, 4.530076, 5.530076, 
    6.530076, 7.530076, 8.530076, 9.530076, 10.53008, 11.53008, 12.53008, 
    13.53008, 14.53008, 15.53008, 16.53008, 17.53008, 18.53008, 19.53008, 
    20.53008, 21.53008, 22.53008, 23.53008, 24.53008, 25.53008, 26.53008, 
    27.53008, 28.53008, 29.53008, 30.53008, 31.53008, 32.53008, 33.53008, 
    34.53008, 35.53008, 36.53008,
  78.00441, 79.00162, 81.99559, 83.99119, 85.98682, 87.98249, 89.97823, 
    91.97403, 93.96992, 95.96591, 97.96202, 99.95825, 101.9546, 103.9512, 
    105.9479, 107.9448, 109.9418, 111.9391, 113.9366, 115.9344, 117.9323, 
    119.9306, 121.9291, 123.9278, 125.9268, 127.9261, 129.9257, 131.9256, 
    133.9257, 135.9261, 137.9268, 139.9278, 141.9291, 143.9306, 145.9324, 
    147.9345, 149.9368, 151.9393, 153.9421, 155.945, 157.9482, 159.9514, 
    161.9549, 163.9585, 165.9622, 167.966, 169.9699, 171.9739, 173.9778, 
    175.9818, 177.9858, 179.9897, -178.0064, -176.0026, -173.9988, -171.9952, 
    -169.9917, -167.9884, -165.9852, -163.9823, -161.9794, -159.9769, 
    -157.9745, -155.9723, -153.9704, -151.9687, -149.9673, -147.9661, 
    -145.9651, -143.9644, -141.964, -139.9638, -137.9639, -135.9642, 
    -133.9647, -131.9655, -129.9665, -127.9677, -125.9691, -123.9707, 
    -121.9725, -119.9745, -117.9766, -115.9788, -113.9812, -111.9837, 
    -109.9862, -107.9889, -105.9916, -103.9944, -101.9972, -100, -98.00282, 
    -96.00562, -94.00839, -92.01112, -90.01377, -88.01635, -86.01883, 
    -84.02119, -82.02344, -80.02554, -78.02749, -76.02927, -74.03087, 
    -72.03228, -70.03349, -68.03448, -66.03526, -64.0358, -62.03611, 
    -60.03617, -58.03599, -56.03556, -54.03487, -52.03393, -50.03274, 
    -48.0313, -46.02962, -44.02769, -42.02554, -40.02316, -38.02056, 
    -36.01775, -34.01476, -32.01159, -30.00825, -28.00477, -26.00115, 
    -23.99743, -21.99362, -19.98973, -17.98579, -15.98182, -13.97783, 
    -11.97386, -9.969924, -8.2199, -6.7199, -5.469924, -4.469924, -3.469924, 
    -2.469924, -1.469924, -0.4699244, 0.5300756, 1.530076, 2.530076, 
    3.530076, 4.530076, 5.530076, 6.530076, 7.530076, 8.530076, 9.530076, 
    10.53008, 11.53008, 12.53008, 13.53008, 14.53008, 15.53008, 16.53008, 
    17.53008, 18.53008, 19.53008, 20.53008, 21.53008, 22.53008, 23.53008, 
    24.53008, 25.53008, 26.53008, 27.53008, 28.53008, 29.53008, 30.53008, 
    31.53008, 32.53008, 33.53008, 34.53008, 35.53008, 36.53008,
  78.00661, 79.00162, 81.99339, 83.98679, 85.98023, 87.97374, 89.96733, 
    91.96102, 93.95483, 95.94878, 97.9429, 99.93721, 101.9317, 103.9264, 
    105.9214, 107.9167, 109.9122, 111.908, 113.9042, 115.9007, 117.8975, 
    119.8947, 121.8923, 123.8903, 125.8888, 127.8876, 129.8868, 131.8865, 
    133.8867, 135.8872, 137.8882, 139.8896, 141.8915, 143.8938, 145.8965, 
    147.8996, 149.903, 151.9068, 153.911, 155.9155, 157.9203, 159.9254, 
    161.9307, 163.9362, 165.9419, 167.9478, 169.9537, 171.9598, 173.9659, 
    175.9721, 177.9782, 179.9843, -178.0097, -176.0038, -173.998, -171.9925, 
    -169.9871, -167.9819, -165.977, -163.9724, -161.9681, -159.9641, 
    -157.9604, -155.9571, -153.9541, -151.9515, -149.9493, -147.9475, 
    -145.9461, -143.9451, -141.9444, -139.9442, -137.9443, -135.9448, 
    -133.9456, -131.9468, -129.9484, -127.9503, -125.9525, -123.9549, 
    -121.9577, -119.9607, -117.9639, -115.9674, -113.9711, -111.9749, 
    -109.9788, -107.9829, -105.9871, -103.9914, -101.9957, -100, -98.00433, 
    -96.00864, -94.01289, -92.01708, -90.02116, -88.02513, -86.02895, 
    -84.0326, -82.03606, -80.0393, -78.04231, -76.04507, -74.04755, 
    -72.04974, -70.05161, -68.05316, -66.05437, -64.05524, -62.05573, 
    -60.05585, -58.05559, -56.05495, -54.05391, -52.05248, -50.05066, 
    -48.04846, -46.04588, -44.04292, -42.03959, -40.03592, -38.03191, 
    -36.02759, -34.02296, -32.01806, -30.01291, -28.00753, -26.00195, 
    -23.99619, -21.9903, -19.98429, -17.9782, -15.97207, -13.96593, -11.9598, 
    -9.953736, -8.21, -6.7154, -5.469924, -4.469924, -3.469924, -2.469924, 
    -1.469924, -0.4699244, 0.5300756, 1.530076, 2.530076, 3.530076, 4.530076, 
    5.530076, 6.530076, 7.530076, 8.530076, 9.530076, 10.53008, 11.53008, 
    12.53008, 13.53008, 14.53008, 15.53008, 16.53008, 17.53008, 18.53008, 
    19.53008, 20.53008, 21.53008, 22.53008, 23.53008, 24.53008, 25.53008, 
    26.53008, 27.53008, 28.53008, 29.53008, 30.53008, 31.53008, 32.53008, 
    33.53008, 34.53008, 35.53008, 36.53008,
  78.00945, 79.00162, 81.99055, 83.98112, 85.97176, 87.96246, 89.95328, 
    91.94423, 93.93535, 95.92665, 97.91818, 99.90995, 101.902, 103.8944, 
    105.8871, 107.8801, 109.8736, 111.8674, 113.8618, 115.8566, 117.8519, 
    119.8477, 121.8441, 123.8411, 125.8386, 127.8368, 129.8355, 131.8349, 
    133.835, 135.8356, 137.837, 139.8389, 141.8415, 143.8447, 145.8485, 
    147.853, 149.8579, 151.8635, 153.8695, 155.8761, 157.883, 159.8904, 
    161.8982, 163.9063, 165.9146, 167.9232, 169.9321, 171.941, 173.95, 
    175.9591, 177.9681, 179.9771, -178.0141, -176.0054, -173.9969, -171.9886, 
    -169.9807, -167.9731, -165.9658, -163.959, -161.9527, -159.9467, 
    -157.9413, -155.9364, -153.9321, -151.9283, -149.9251, -147.9224, 
    -145.9204, -143.9189, -141.918, -139.9176, -137.9178, -135.9186, 
    -133.9199, -131.9217, -129.924, -127.9268, -125.93, -123.9337, -121.9378, 
    -119.9422, -117.947, -115.9521, -113.9575, -111.9631, -109.9689, 
    -107.9749, -105.9811, -103.9873, -101.9936, -100, -98.00636, -96.01268, 
    -94.01893, -92.02507, -90.03107, -88.0369, -86.04252, -84.04789, 
    -82.05298, -80.05776, -78.06221, -76.06628, -74.06995, -72.0732, 
    -70.07599, -68.07831, -66.08012, -64.08142, -62.08218, -60.0824, 
    -58.08205, -56.08113, -54.07964, -52.07756, -50.07491, -48.07168, 
    -46.06789, -44.06355, -42.05866, -40.05326, -38.04735, -36.04098, 
    -34.03416, -32.02693, -30.01932, -28.01138, -26.00314, -23.99464, 
    -21.98594, -19.97708, -17.9681, -15.95905, -13.95, -11.94098, -9.932048, 
    -8.199539, -6.71315, -5.467674, -4.469924, -3.469924, -2.469924, 
    -1.469924, -0.4699244, 0.5300756, 1.530076, 2.530076, 3.530076, 4.530076, 
    5.530076, 6.530076, 7.530076, 8.530076, 9.530076, 10.53008, 11.53008, 
    12.53008, 13.53008, 14.53008, 15.53008, 16.53008, 17.53008, 18.53008, 
    19.53008, 20.53008, 21.53008, 22.53008, 23.53008, 24.53008, 25.53008, 
    26.53008, 27.53008, 28.53008, 29.53008, 30.53008, 31.53008, 32.53008, 
    33.53008, 34.53008, 35.53008, 36.53008,
  78.01298, 80, 81.98702, 83.97408, 85.9612, 87.94843, 89.93578, 91.92331, 
    93.91103, 95.89901, 97.88726, 99.87583, 101.8648, 103.8541, 105.8439, 
    107.8341, 109.8249, 111.8162, 113.8081, 115.8007, 117.794, 119.788, 
    121.7827, 123.7782, 125.7746, 127.7718, 129.7698, 131.7688, 133.7686, 
    135.7693, 137.771, 139.7736, 141.777, 143.7814, 145.7866, 147.7927, 
    149.7996, 151.8073, 153.8158, 155.8249, 157.8347, 159.8451, 161.856, 
    163.8674, 165.8793, 167.8914, 169.9039, 171.9166, 173.9294, 175.9422, 
    177.9551, 179.9678, -178.0196, -176.0072, -173.9951, -171.9834, 
    -169.9721, -167.9613, -165.951, -163.9413, -161.9323, -159.9239, 
    -157.9162, -155.9093, -153.9032, -151.8978, -149.8933, -147.8896, 
    -145.8867, -143.8846, -141.8833, -139.8829, -137.8832, -135.8844, 
    -133.8863, -131.8889, -129.8922, -127.8962, -125.9009, -123.9061, 
    -121.9119, -119.9182, -117.925, -115.9322, -113.9399, -111.9478, 
    -109.9561, -107.9646, -105.9732, -103.9821, -101.991, -100, -98.00899, 
    -96.01792, -94.02676, -92.03545, -90.04395, -88.05219, -86.06014, 
    -84.06776, -82.07499, -80.08178, -78.0881, -76.0939, -74.09914, 
    -72.10378, -70.10777, -68.11111, -66.11373, -64.11562, -62.11675, 
    -60.11711, -58.11666, -56.11541, -54.11333, -52.11043, -50.1067, 
    -48.10216, -46.09681, -44.09066, -42.08375, -40.07609, -38.06771, 
    -36.05866, -34.04897, -32.0387, -30.02789, -28.01659, -26.00488, 
    -23.9928, -21.98042, -19.96782, -17.95506, -15.94222, -13.92936, 
    -11.91656, -9.903902, -8.029911, -6.316759, -4.687521, -4.469924, 
    -3.469924, -2.469924, -1.469924, -0.4699244, 0.5300756, 1.530076, 
    2.530076, 3.530076, 4.530076, 5.530076, 6.530076, 7.530076, 8.530076, 
    9.530076, 10.53008, 11.53008, 12.53008, 13.53008, 14.53008, 15.53008, 
    16.53008, 17.53008, 18.53008, 19.53008, 20.53008, 21.53008, 22.53008, 
    23.53008, 24.53008, 25.53008, 26.53008, 27.53008, 28.53008, 29.53008, 
    30.53008, 31.53008, 32.53008, 33.53008, 34.53008, 35.53008, 80,
  78.01723, 80, 81.98277, 83.96557, 85.94845, 87.93144, 89.9146, 91.89796, 
    93.88155, 95.86545, 97.84968, 99.8343, 101.8194, 103.8049, 105.791, 
    107.7777, 109.7651, 111.7532, 113.7421, 115.7318, 117.7225, 119.714, 
    121.7066, 123.7003, 125.695, 127.6909, 129.6879, 131.6862, 133.6856, 
    135.6864, 137.6883, 139.6916, 141.6961, 143.7018, 145.7087, 147.7168, 
    149.7261, 151.7365, 153.7479, 155.7603, 157.7736, 159.7878, 161.8027, 
    163.8183, 165.8345, 167.8512, 169.8683, 171.8857, 173.9033, 175.921, 
    177.9387, 179.9563, -178.0264, -176.0093, -173.9927, -171.9765, -169.961, 
    -167.946, -165.9319, -163.9186, -161.9061, -159.8946, -157.8841, 
    -155.8746, -153.8661, -151.8588, -149.8526, -147.8476, -145.8436, 
    -143.8409, -141.8392, -139.8387, -137.8392, -135.8408, -133.8435, 
    -131.8472, -129.8518, -127.8574, -125.8638, -123.8711, -121.8791, 
    -119.8878, -117.8971, -115.9071, -113.9175, -111.9285, -109.9398, 
    -107.9514, -105.9633, -103.9754, -101.9877, -100, -98.01231, -96.02455, 
    -94.03667, -92.04858, -90.06023, -88.07155, -86.08247, -84.09293, 
    -82.10287, -80.11223, -78.12094, -76.12894, -74.13619, -72.14262, 
    -70.14817, -68.15282, -66.15649, -64.15916, -62.16079, -60.16135, 
    -58.16081, -56.15916, -54.15637, -52.15244, -50.14737, -48.14117, 
    -46.13384, -44.12542, -42.11593, -40.1054, -38.09389, -36.08144, 
    -34.0681, -32.05395, -30.03905, -28.02349, -26.00734, -23.99069, 
    -21.97364, -19.95628, -17.93871, -15.92102, -13.90333, -11.88573, 
    -9.868335, -7.851233, -5.83453, -3.818324, -4.469924, -3.469924, 
    -2.469924, -1.469924, -0.4699244, 0.5300756, 1.530076, 2.530076, 
    3.530076, 4.530076, 5.530076, 6.530076, 7.530076, 8.530076, 9.530076, 
    10.53008, 11.53008, 12.53008, 13.53008, 14.53008, 15.53008, 16.53008, 
    17.53008, 18.53008, 19.53008, 20.53008, 21.53008, 22.53008, 23.53008, 
    24.53008, 25.53008, 26.53008, 27.53008, 28.53008, 29.53008, 30.53008, 
    31.53008, 32.53008, 33.53008, 34.53008, 35.53008, 80,
  78.02225, 80, 81.97775, 83.95554, 85.9334, 87.91141, 89.88958, 91.86798, 
    93.84666, 95.82566, 97.80506, 99.78491, 101.7653, 103.7462, 105.7279, 
    107.7102, 109.6934, 111.6775, 113.6626, 115.6488, 117.636, 119.6245, 
    121.6144, 123.6055, 125.5982, 127.5923, 129.588, 131.5852, 133.5841, 
    135.5847, 137.5869, 139.5909, 141.5965, 143.6038, 145.6127, 147.6233, 
    149.6354, 151.649, 153.664, 155.6804, 157.6981, 159.7169, 161.7368, 
    163.7576, 165.7792, 167.8015, 169.8244, 171.8477, 173.8712, 175.8949, 
    177.9187, 179.9422, -178.0345, -176.0116, -173.9892, -171.9676, 
    -169.9467, -167.9267, -165.9077, -163.8898, -161.8731, -159.8577, 
    -157.8436, -155.831, -153.8197, -151.81, -149.8017, -147.795, -145.7898, 
    -143.7862, -141.7841, -139.7834, -137.7843, -135.7866, -133.7903, 
    -131.7953, -129.8016, -127.8091, -125.8178, -123.8275, -121.8383, 
    -119.85, -117.8625, -115.8759, -113.8899, -111.9045, -109.9196, 
    -107.9352, -105.9511, -103.9672, -101.9836, -100, -98.01643, -96.03276, 
    -94.04893, -92.06483, -90.0804, -88.09552, -86.11013, -84.12414, 
    -82.13746, -80.15001, -78.16171, -76.17248, -74.18224, -72.19091, 
    -70.19843, -68.20473, -66.20975, -64.21342, -62.21571, -60.21656, 
    -58.21594, -56.21381, -54.21017, -52.20499, -50.19828, -48.19003, 
    -46.18028, -44.16904, -42.15636, -40.14227, -38.12685, -36.11017, 
    -34.09229, -32.07331, -30.05332, -28.03243, -26.01076, -23.98842, 
    -21.96553, -19.94224, -17.91866, -15.89495, -13.87124, -11.84767, 
    -9.824379, -7.80151, -5.779197, -3.757573, -1.736766, 0.2831027, 
    0.3831027, 0.4831027, -0.4699244, 0.5300756, 1.530076, 2.530076, 
    3.530076, 4.530076, 5.530076, 6.530076, 7.530076, 8.530076, 9.530076, 
    10.53008, 11.53008, 12.53008, 13.53008, 14.53008, 15.53008, 16.53008, 
    17.53008, 18.53008, 19.53008, 20.53008, 21.53008, 22.53008, 23.53008, 
    24.53008, 25.53008, 26.53008, 27.53008, 28.53008, 29.53008, 30.53008, 
    31.53008, 32.53008, 33.53008, 34.53008, 35.53008, 80,
  78.02805, 80, 81.97195, 83.94395, 85.91604, 87.88825, 89.86065, 91.83327, 
    93.80618, 95.77945, 97.75314, 99.72734, 101.7021, 103.6776, 105.6538, 
    107.631, 109.609, 111.5882, 113.5686, 115.5503, 117.5335, 119.5182, 
    121.5045, 123.4926, 125.4825, 127.4743, 129.4682, 131.4641, 133.4621, 
    135.4624, 137.4648, 139.4694, 141.4763, 143.4854, 145.4966, 147.51, 
    149.5255, 151.543, 153.5624, 155.5836, 157.6064, 159.6309, 161.6567, 
    163.6838, 165.712, 167.7412, 169.7711, 171.8016, 173.8324, 175.8635, 
    177.8946, 179.9255, -178.0439, -176.0139, -173.9846, -171.9562, 
    -169.9288, -167.9025, -165.8776, -163.8542, -161.8324, -159.8122, 
    -157.7938, -155.7772, -153.7625, -151.7498, -149.7391, -147.7304, 
    -145.7238, -143.7191, -141.7165, -139.7158, -137.717, -135.7202, 
    -133.7251, -131.7318, -129.7402, -127.7501, -125.7616, -123.7744, 
    -121.7886, -119.804, -117.8204, -115.8379, -113.8562, -111.8753, 
    -109.8951, -107.9154, -105.9362, -103.9573, -101.9786, -100, -98.02142, 
    -96.04274, -94.06384, -92.0846, -90.10492, -88.12469, -86.1438, 
    -84.16213, -82.17958, -80.19604, -78.21141, -76.22557, -74.23843, 
    -72.24988, -70.25983, -68.2682, -66.27489, -64.27985, -62.28297, 
    -60.28422, -58.28354, -56.28089, -54.27624, -52.26957, -50.26088, 
    -48.25017, -46.23746, -44.22281, -42.20624, -40.18782, -38.16764, 
    -36.14579, -34.12235, -32.09747, -30.07125, -28.04384, -26.01541, 
    -23.98609, -21.95606, -19.9255, -17.89458, -15.8635, -13.83243, 
    -11.80156, -9.771079, -7.741177, -5.71203, -3.683817, -1.656705, 
    0.3691426, 0.4691426, 0.5691426, 0.6691426, 0.5300756, 1.530076, 
    2.530076, 3.530076, 4.530076, 5.530076, 6.530076, 7.530076, 8.530076, 
    9.530076, 10.53008, 11.53008, 12.53008, 13.53008, 14.53008, 15.53008, 
    16.53008, 17.53008, 18.53008, 19.53008, 20.53008, 21.53008, 22.53008, 
    23.53008, 24.53008, 25.53008, 26.53008, 27.53008, 28.53008, 29.53008, 
    30.53008, 31.53008, 32.53008, 33.53008, 34.53008, 35.53008, 80,
  78.0346, 80, 81.9654, 83.93084, 85.89635, 87.86198, 89.82776, 91.79376, 
    93.76005, 95.72668, 97.69375, 99.66135, 101.6296, 103.5986, 105.5684, 
    107.5393, 109.5113, 111.4846, 113.4593, 115.4356, 117.4137, 119.3936, 
    121.3756, 123.3598, 125.3463, 127.3353, 129.3267, 131.3209, 133.3177, 
    135.3174, 137.3198, 139.3252, 141.3334, 143.3445, 145.3584, 147.3751, 
    149.3945, 151.4165, 153.441, 155.4678, 157.4969, 159.528, 161.561, 
    163.5957, 165.6318, 167.6691, 169.7075, 171.7466, 173.7863, 175.8262, 
    177.8662, 179.9059, -178.0547, -176.0161, -173.9784, -171.9418, 
    -169.9065, -167.8728, -165.8408, -163.8107, -161.7826, -159.7567, 
    -157.7331, -155.7119, -153.6932, -151.6769, -149.6633, -147.6523, 
    -145.6439, -143.6381, -141.6348, -139.6341, -137.6359, -135.6401, 
    -133.6466, -131.6554, -129.6663, -127.6792, -125.6941, -123.7107, 
    -121.7289, -119.7487, -117.7699, -115.7923, -113.8159, -111.8404, 
    -109.8657, -107.8917, -105.9183, -103.9453, -101.9726, -100, -98.02741, 
    -96.05468, -94.08167, -92.10826, -90.13428, -88.15962, -86.18413, 
    -84.20766, -82.23009, -80.25127, -78.27106, -76.28933, -74.30595, 
    -72.32078, -70.3337, -68.3446, -66.35337, -64.35989, -62.36409, 
    -60.36587, -58.36518, -56.36194, -54.35613, -52.34771, -50.33669, 
    -48.32305, -46.30684, -44.28809, -42.26688, -40.24326, -38.21736, 
    -36.18929, -34.15917, -32.12717, -30.09345, -28.0582, -26.0216, 
    -23.98388, -21.94525, -19.90593, -17.86616, -15.82619, -13.78626, 
    -11.74661, -9.707494, -7.669143, -5.631798, -3.595689, -1.561035, 
    0.4719526, 0.5719526, 0.6719526, 0.7719526, 0.8719526, 1.530076, 
    2.530076, 3.530076, 4.530076, 5.530076, 6.530076, 7.530076, 8.530076, 
    9.530076, 10.53008, 11.53008, 12.53008, 13.53008, 14.53008, 15.53008, 
    16.53008, 17.53008, 18.53008, 19.53008, 20.53008, 21.53008, 22.53008, 
    23.53008, 24.53008, 25.53008, 26.53008, 27.53008, 28.53008, 29.53008, 
    30.53008, 31.53008, 32.53008, 33.53008, 34.53008, 35.53008, 80,
  78.04191, 80, 81.95809, 83.91621, 85.87437, 87.83261, 89.79097, 91.74949, 
    93.70824, 95.6673, 97.62677, 99.58675, 101.5474, 103.5088, 105.4712, 
    107.4346, 109.3994, 111.3657, 113.3336, 115.3035, 117.2754, 119.2497, 
    121.2264, 123.2058, 125.1881, 127.1734, 129.1619, 131.1537, 133.1489, 
    135.1477, 137.1501, 139.1561, 141.1657, 143.179, 145.1959, 147.2163, 
    149.2402, 151.2675, 153.298, 155.3315, 157.3679, 159.4069, 161.4483, 
    163.4918, 165.5373, 167.5843, 169.6327, 171.6821, 173.7321, 175.7826, 
    177.8331, 179.8834, -178.0668, -176.018, -173.9703, -171.924, -169.8794, 
    -167.8367, -165.7963, -163.7583, -161.7228, -159.6901, -157.6604, 
    -155.6337, -153.6101, -151.5898, -149.5727, -147.5589, -145.5485, 
    -143.5414, -141.5375, -139.5369, -137.5394, -135.5449, -133.5534, 
    -131.5646, -129.5786, -127.5951, -125.614, -123.6351, -121.6583, 
    -119.6834, -117.7101, -115.7385, -113.7682, -111.7991, -109.831, 
    -107.8638, -105.8973, -103.9312, -101.9655, -100, -98.03447, -96.06878, 
    -94.10274, -92.1362, -90.16898, -88.2009, -86.23181, -84.26152, 
    -82.28986, -80.31664, -78.34171, -76.36489, -74.386, -72.40489, 
    -70.42139, -68.43536, -66.44664, -64.45511, -62.46064, -60.46312, 
    -58.46247, -56.45861, -54.45148, -52.44105, -50.4273, -48.41024, 
    -46.38991, -44.36634, -42.33963, -40.30988, -38.2772, -36.24175, 
    -34.20371, -32.16326, -30.12062, -28.07604, -26.02975, -23.98202, 
    -21.93315, -19.88342, -17.83313, -15.78261, -13.73215, -11.68207, 
    -9.632695, -7.584328, -5.537273, -3.491823, -1.448261, 0.5931457, 
    0.6931457, 0.7931457, 0.8931457, 0.9931456, 1.530076, 2.530076, 3.530076, 
    4.530076, 5.530076, 6.530076, 7.530076, 8.530076, 9.530076, 10.53008, 
    11.53008, 12.53008, 13.53008, 14.53008, 15.53008, 16.53008, 17.53008, 
    18.53008, 19.53008, 20.53008, 21.53008, 22.53008, 23.53008, 24.53008, 
    25.53008, 26.53008, 27.53008, 28.53008, 29.53008, 30.53008, 31.53008, 
    32.53008, 33.53008, 34.53008, 35.53008, 80,
  78.04994, 80, 81.95006, 83.90012, 85.85017, 87.80024, 89.75034, 91.7005, 
    93.65079, 95.60131, 97.55215, 99.50343, 101.4553, 103.408, 105.3617, 
    107.3165, 109.2729, 111.2308, 113.1908, 115.1529, 117.1176, 119.085, 
    121.0554, 123.029, 125.0061, 126.987, 128.9718, 130.9607, 132.9538, 
    134.9514, 136.9534, 138.9599, 140.9711, 142.9868, 145.007, 147.0317, 
    149.0608, 151.0941, 153.1315, 155.1727, 157.2175, 159.2657, 161.3169, 
    163.3708, 165.4272, 167.4857, 169.5458, 171.6072, 173.6695, 175.7323, 
    177.7953, 179.8579, -178.0801, -176.0192, -173.9597, -171.902, -169.8465, 
    -167.7934, -165.743, -163.6957, -161.6516, -159.611, -157.574, -155.5409, 
    -153.5117, -151.4866, -149.4656, -147.4487, -145.436, -143.4274, 
    -141.4229, -139.4224, -137.4258, -135.4329, -133.4438, -131.4581, 
    -129.4757, -127.4965, -125.5202, -123.5466, -121.5756, -119.6069, 
    -117.6403, -115.6755, -113.7125, -111.7509, -109.7905, -107.8312, 
    -105.8727, -103.9148, -101.9573, -100, -98.04272, -96.08522, -94.12733, 
    -92.16882, -90.20949, -88.24912, -86.28753, -84.32447, -82.35975, 
    -80.39314, -78.42443, -76.4534, -74.47984, -72.50355, -70.52431, 
    -68.54194, -66.55624, -64.56706, -62.57424, -60.57763, -58.57711, 
    -56.57259, -54.564, -52.55127, -50.5344, -48.51339, -46.48826, -44.45909, 
    -42.42597, -40.38903, -38.34843, -36.30434, -34.257, -32.20664, 
    -30.15353, -28.09797, -26.04029, -23.98081, -21.91989, -19.85792, 
    -17.79527, -15.73233, -13.6695, -11.60718, -9.545772, -7.485659, 
    -5.427228, -3.37085, -1.316878, 0.7343502, 0.8343502, 0.9343502, 1.03435, 
    1.13435, 1.530076, 2.530076, 3.530076, 4.530076, 5.530076, 6.530076, 
    7.530076, 8.530076, 9.530076, 10.53008, 11.53008, 12.53008, 13.53008, 
    14.53008, 15.53008, 16.53008, 17.53008, 18.53008, 19.53008, 20.53008, 
    21.53008, 22.53008, 23.53008, 24.53008, 25.53008, 26.53008, 27.53008, 
    28.53008, 29.53008, 30.53008, 31.53008, 32.53008, 33.53008, 34.53008, 
    35.53008, 80,
  78.05866, 80, 81.94134, 83.88263, 85.82384, 87.76496, 89.70597, 91.64689, 
    93.58778, 95.52872, 97.46984, 99.41127, 101.3532, 103.2959, 105.2395, 
    107.1844, 109.1309, 111.0793, 113.0298, 114.9829, 116.939, 118.8982, 
    120.8611, 122.8278, 124.7988, 126.7743, 128.7546, 130.7399, 132.7304, 
    134.7262, 136.7276, 138.7346, 140.7473, 142.7656, 144.7896, 146.8191, 
    148.854, 150.8942, 152.9394, 154.9895, 157.044, 159.1028, 161.1654, 
    163.2314, 165.3004, 167.3721, 169.4458, 171.5212, 173.5978, 175.675, 
    177.7524, 179.8294, -178.0943, -176.0194, -173.9462, -171.8753, -169.807, 
    -167.7417, -165.6798, -163.6217, -161.5676, -159.5178, -157.4725, 
    -155.432, -153.3964, -151.3658, -149.3402, -147.3198, -145.3045, 
    -143.2943, -141.2891, -139.2889, -137.2934, -135.3026, -133.3162, 
    -131.3342, -129.3561, -127.3819, -125.4113, -123.4439, -121.4797, 
    -119.5182, -117.5593, -115.6027, -113.648, -111.6951, -109.7437, 
    -107.7935, -105.8443, -103.8958, -101.9478, -100, -98.05223, -96.10423, 
    -94.15573, -92.2065, -90.25631, -88.30489, -86.35197, -84.39732, 
    -82.44067, -80.48176, -78.5203, -76.55605, -74.58874, -72.6181, 
    -70.64388, -68.66585, -66.68376, -64.69741, -62.70659, -60.71112, 
    -58.71087, -56.70568, -54.69547, -52.68017, -50.65975, -48.63421, 
    -46.60359, -44.56797, -42.52746, -40.48221, -38.43242, -36.37832, 
    -34.32018, -32.2583, -30.19302, -28.1247, -26.05375, -23.98059, 
    -21.90566, -19.82943, -17.75238, -15.675, -13.59778, -11.52122, 
    -9.445818, -7.372064, -5.300432, -3.231384, -1.165361, 0.89722, 0.99722, 
    1.09722, 1.19722, 1.29722, 1.530076, 2.530076, 3.530076, 4.530076, 
    5.530076, 6.530076, 7.530076, 8.530076, 9.530076, 10.53008, 11.53008, 
    12.53008, 13.53008, 14.53008, 15.53008, 16.53008, 17.53008, 18.53008, 
    19.53008, 20.53008, 21.53008, 22.53008, 23.53008, 24.53008, 25.53008, 
    26.53008, 27.53008, 28.53008, 29.53008, 30.53008, 31.53008, 32.53008, 
    33.53008, 34.53008, 35.53008, 80,
  78.06804, 80, 81.93196, 83.86382, 85.79549, 87.7269, 89.658, 91.58878, 
    93.51928, 95.44958, 97.37981, 99.31014, 101.2408, 103.1721, 105.1043, 
    107.0378, 108.9729, 110.91, 112.8497, 114.7923, 116.7383, 118.688, 
    120.642, 122.6006, 124.5643, 126.5334, 128.5083, 130.4892, 132.4764, 
    134.4702, 136.4706, 138.4779, 140.4922, 142.5133, 144.5414, 146.5762, 
    148.6177, 150.6657, 152.7199, 154.78, 156.8457, 158.9165, 160.9922, 
    163.072, 165.1556, 167.2425, 169.3319, 171.4235, 173.5164, 175.6103, 
    177.7043, 179.798, -178.1093, -176.0182, -173.9292, -171.843, -169.7599, 
    -167.6806, -165.6055, -163.5349, -161.4693, -159.409, -157.3542, 
    -155.3053, -153.2623, -151.2254, -149.1948, -147.1704, -145.1522, 
    -143.1403, -141.1344, -139.1346, -137.1405, -135.1521, -133.1692, 
    -131.1913, -129.2184, -127.25, -125.286, -123.3259, -121.3695, -119.4165, 
    -117.4664, -115.5191, -113.5741, -111.6312, -109.69, -107.7503, 
    -105.8117, -103.874, -101.9369, -100, -98.06313, -96.12598, -94.18826, 
    -92.24968, -90.30995, -88.36878, -86.42587, -84.4809, -82.53355, 
    -80.58351, -78.63046, -76.67406, -74.714, -72.74995, -70.78161, 
    -68.80867, -66.83083, -64.84785, -62.85946, -60.86543, -58.86558, 
    -56.85974, -54.84779, -52.82963, -50.80523, -48.77458, -46.73771, 
    -44.69473, -42.64576, -40.591, -38.53067, -36.46507, -34.3945, -32.31936, 
    -30.24005, -28.15702, -26.07076, -23.98181, -21.8907, -19.79801, 
    -17.70433, -15.61027, -13.51645, -11.42346, -9.331932, -7.24246, 
    -5.155632, -3.072016, -0.9921508, 1.083451, 3.154314, 5.220001, 7.280117, 
    9.334314, 11.38229, 13.4238, 15.45865, 17.48669, 19.50784, 21.52206, 
    23.52937, 25.52984, 27.52361, 29.51083, 31.49174, 33.46659, 35.43569, 
    37.39937, 39.35801, 41.31199, 17.53008, 18.53008, 19.53008, 20.53008, 
    21.53008, 22.53008, 23.53008, 24.53008, 25.53008, 26.53008, 27.53008, 
    28.53008, 29.53008, 30.53008, 31.53008, 32.53008, 33.53008, 34.53008, 
    35.53008, 80,
  78.07802, 80, 81.92198, 83.84379, 85.76524, 87.68619, 89.60654, 91.52627, 
    93.44534, 95.36387, 97.28197, 99.19987, 101.1178, 103.0362, 104.9554, 
    106.8758, 108.7979, 110.7222, 112.6493, 114.5798, 116.5141, 118.4528, 
    120.3964, 122.3456, 124.3007, 126.2623, 128.2308, 130.2065, 132.1897, 
    134.1808, 136.1801, 138.1875, 140.2033, 142.2275, 144.26, 146.3008, 
    148.3497, 150.4064, 152.4707, 154.5423, 156.6206, 158.7052, 160.7956, 
    162.8913, 164.9915, 167.0957, 169.2032, 171.3132, 173.425, 175.5379, 
    177.651, 179.7638, -178.1247, -176.015, -173.908, -171.8042, -169.7043, 
    -167.609, -165.5187, -163.4339, -161.3552, -159.2829, -157.2173, 
    -155.1588, -153.1075, -151.0636, -149.0272, -146.9983, -144.9771, 
    -142.9632, -140.9568, -138.9576, -136.9653, -134.9798, -133.0008, 
    -131.028, -129.061, -127.0994, -125.143, -123.1913, -121.244, -119.3005, 
    -117.3607, -115.424, -113.4901, -111.5585, -109.6291, -107.7013, 
    -105.7748, -103.8493, -101.9245, -100, -98.07551, -96.15068, -94.2252, 
    -92.29874, -90.37094, -88.44146, -86.50994, -84.57602, -82.63932, 
    -80.69946, -78.75604, -76.80868, -74.85699, -72.90056, -70.93903, 
    -68.97202, -66.99918, -65.02016, -63.03468, -61.04244, -59.0432, 
    -57.03675, -55.02295, -53.00166, -50.97283, -48.93645, -46.89256, 
    -44.84125, -42.7827, -40.71713, -38.64481, -36.56608, -34.48134, 
    -32.39104, -30.29568, -28.1958, -26.09203, -23.98497, -21.87532, 
    -19.76376, -17.65103, -15.53786, -13.425, -11.3132, -9.2032, -7.095745, 
    -4.991544, -2.891288, -0.7956332, 1.294801, 3.37944, 5.457756, 7.529276, 
    9.593583, 11.65032, 13.6992, 15.73998, 17.77251, 19.79669, 21.81249, 
    23.81994, 25.81915, 27.81028, 29.79355, 31.76925, 33.73769, 35.69926, 
    37.6544, 39.60356, 41.54723, 17.53008, 18.53008, 19.53008, 20.53008, 
    21.53008, 22.53008, 23.53008, 24.53008, 25.53008, 26.53008, 27.53008, 
    28.53008, 29.53008, 30.53008, 31.53008, 32.53008, 33.53008, 34.53008, 
    35.53008, 80,
  78.08855, 80, 81.91145, 83.8226, 85.73318, 87.64295, 89.55174, 91.45944, 
    93.36603, 95.27157, 97.17621, 99.08022, 100.9839, 102.8877, 104.7921, 
    106.6977, 108.605, 110.5147, 112.4274, 114.3439, 116.2648, 118.1908, 
    120.1226, 122.0608, 124.0061, 125.9589, 127.9199, 129.8894, 131.868, 
    133.8559, 135.8535, 137.8609, 139.8783, 141.9057, 143.9431, 145.9905, 
    148.0475, 150.1141, 152.1897, 154.2741, 156.3667, 158.4669, 160.5741, 
    162.6877, 164.8068, 166.9308, 169.0587, 171.1897, 173.3229, 175.4575, 
    177.5924, 179.7269, -178.1401, -176.0093, -173.8816, -171.7579, 
    -169.6389, -167.5253, -165.4178, -163.317, -161.2234, -159.1375, 
    -157.0598, -154.9904, -152.9298, -150.8781, -148.8353, -146.8016, 
    -144.7769, -142.7612, -140.7542, -138.7558, -136.7658, -134.7838, 
    -132.8094, -130.8424, -128.8822, -126.9286, -124.9809, -123.0388, 
    -121.1018, -119.1693, -117.2411, -115.3164, -113.3951, -111.4765, 
    -109.5602, -107.6459, -105.7331, -103.8214, -101.9105, -100, -98.08947, 
    -96.17856, -94.26691, -92.35411, -90.43979, -88.52354, -86.60493, 
    -84.68356, -82.75895, -80.83067, -78.89825, -76.96121, -75.0191, 
    -73.07143, -71.11776, -69.15762, -67.19057, -65.21623, -63.23421, 
    -61.24416, -59.24578, -57.23882, -55.22307, -53.19839, -51.16469, 
    -49.12194, -47.0702, -45.00957, -42.94025, -40.86248, -38.77661, 
    -36.68303, -34.58221, -32.4747, -30.3611, -28.24208, -26.11836, -23.9907, 
    -21.85992, -19.72687, -17.59242, -15.45747, -13.32293, -11.1897, 
    -9.058684, -6.930774, -4.806829, -2.68768, -0.5741176, 1.533115, 3.63333, 
    5.725898, 7.810256, 9.885913, 11.95245, 14.00952, 16.05687, 18.0943, 
    20.12173, 22.13911, 24.14652, 26.14408, 28.13201, 30.11058, 32.08014, 
    34.0411, 35.99394, 37.93918, 39.87739, 41.80918, 43.7352, 45.6561, 
    47.57258, 49.48533, 51.39502, 53.30232, 55.20787, 57.11228, 59.01609, 
    60.91979, 62.82379, 64.72843, 66.63397, 68.54056, 70.44826, 72.35705, 
    74.26682, 76.1774, 78.08855, 80,
  78.0996, 80, 81.9004, 83.80035, 85.69945, 87.59732, 89.49368, 91.38837, 
    93.28131, 95.17255, 97.06229, 98.95081, 100.8385, 102.726, 104.6137, 
    106.5025, 108.393, 110.2861, 112.1825, 114.0831, 115.9888, 117.9003, 
    119.8185, 121.7442, 123.6781, 125.6209, 127.5732, 129.5357, 131.5087, 
    133.4928, 135.4883, 137.4955, 139.5145, 141.5453, 143.5881, 145.6427, 
    147.7088, 149.7863, 151.8746, 153.9733, 156.0819, 158.1996, 160.3258, 
    162.4596, 164.6001, 166.7464, 168.8974, 171.0522, 173.2097, 175.3689, 
    177.5285, 179.6876, -178.155, -176.0003, -173.8493, -171.703, -169.5623, 
    -167.4281, -165.3012, -163.1823, -161.072, -158.9709, -156.8795, 
    -154.7981, -152.7271, -150.6666, -148.6169, -146.5779, -144.5496, 
    -142.5318, -140.5245, -138.5273, -136.5399, -134.562, -132.5931, 
    -130.6328, -128.6805, -126.7358, -124.7982, -122.867, -120.9417, 
    -119.0217, -117.1066, -115.1956, -113.2884, -111.3843, -109.4829, 
    -107.5838, -105.6863, -103.7902, -101.8949, -100, -98.10513, -96.20982, 
    -94.31367, -92.41624, -90.51706, -88.61568, -86.71163, -84.80439, 
    -82.89345, -80.97827, -79.05831, -77.13301, -75.20181, -73.26415, 
    -71.31947, -69.36723, -67.40691, -65.43802, -63.46009, -61.47271, 
    -59.47551, -57.46817, -55.45044, -53.42212, -51.38311, -49.33336, 
    -47.27292, -45.20192, -43.12055, -41.02913, -38.92803, -36.81774, 
    -34.69881, -32.57188, -30.43768, -28.29699, -26.15069, -23.9997, 
    -21.84498, -19.68756, -17.5285, -15.36886, -13.20974, -11.05223, 
    -8.897408, -6.746346, -4.600071, -2.459578, -0.3258093, 1.800352, 
    3.918089, 6.026659, 8.1254, 10.21373, 12.29118, 14.35733, 16.4119, 
    18.45468, 20.48556, 22.50453, 24.51167, 26.50716, 28.49127, 30.46432, 
    32.42677, 34.3791, 36.3219, 38.25579, 40.18148, 42.09969, 44.01123, 
    45.91689, 47.81751, 49.71393, 51.60699, 53.49751, 55.38628, 57.27404, 
    59.16148, 61.04919, 62.93771, 64.82745, 66.71869, 68.61163, 70.50632, 
    72.40268, 74.30055, 76.19965, 78.0996, 80,
  78.11111, 80, 81.88889, 83.77714, 85.66414, 87.54938, 89.43243, 91.31305, 
    93.19109, 95.06663, 96.93986, 98.81114, 100.681, 102.5501, 104.4192, 
    106.289, 108.1606, 110.0349, 111.9129, 113.7956, 115.684, 117.5792, 
    119.482, 121.3935, 123.3145, 125.2459, 127.1883, 129.1426, 131.1093, 
    133.0889, 135.0819, 137.0885, 139.109, 141.1436, 143.1922, 145.2547, 
    147.3308, 149.4203, 151.5228, 153.6376, 155.764, 157.9014, 160.0488, 
    162.2052, 164.3698, 166.5412, 168.7183, 170.9, 173.0849, 175.2718, 
    177.4593, 179.6461, -178.1689, -175.9872, -173.8099, -171.6382, 
    -169.4731, -167.3157, -165.167, -163.0277, -160.8988, -158.7807, 
    -156.674, -154.5793, -152.4968, -150.4268, -148.3694, -146.3247, 
    -144.2925, -142.2728, -140.2653, -138.2696, -136.2855, -134.3124, 
    -132.3498, -130.3972, -128.4541, -126.5196, -124.5933, -122.6745, 
    -120.7625, -118.8566, -116.9561, -115.0606, -113.1692, -111.2814, 
    -109.3967, -107.5144, -105.6342, -103.7553, -101.8774, -100, -98.12258, 
    -96.24469, -94.36584, -92.48556, -90.60331, -88.71858, -86.83082, 
    -84.93945, -83.04386, -81.14343, -79.23753, -77.32549, -75.40665, 
    -73.48036, -71.54594, -69.60275, -67.65018, -65.68761, -63.71451, 
    -61.73036, -59.73472, -57.7272, -55.70748, -53.67532, -51.63058, 
    -49.57319, -47.50319, -45.4207, -43.32597, -41.21934, -39.10125, 
    -36.97226, -34.83302, -32.68428, -30.52691, -28.36185, -26.19011, 
    -24.01279, -21.83107, -19.64615, -17.45929, -15.27178, -13.08491, -10.9, 
    -8.718332, -6.541174, -4.369754, -2.205249, -0.04877643, 2.098622, 
    4.235984, 6.362441, 8.47722, 10.57965, 12.66918, 14.74535, 16.80783, 
    18.8564, 20.89095, 22.91149, 24.91813, 26.91109, 28.8907, 30.85738, 
    32.81165, 34.75413, 36.68549, 38.60649, 40.51797, 42.42083, 44.31597, 
    46.2044, 48.08709, 49.96508, 51.83938, 53.71098, 55.58085, 57.44991, 
    59.31899, 61.18885, 63.06015, 64.93337, 66.80891, 68.68695, 70.56757, 
    72.45062, 74.33586, 76.22286, 78.11111, 80,
  78.12305, 80, 81.87695, 83.75301, 85.62733, 87.49919, 89.368, 91.23341, 
    93.09521, 94.95346, 96.80843, 98.66057, 100.5105, 102.3591, 104.2072, 
    106.0559, 107.9062, 109.7595, 111.6168, 113.4794, 115.3484, 117.2252, 
    119.1108, 121.0063, 122.9128, 124.8312, 126.7625, 128.7075, 130.6669, 
    132.6413, 134.6312, 136.6371, 138.6591, 140.6975, 142.7524, 144.8235, 
    146.9107, 149.0135, 151.1316, 153.2641, 155.4105, 157.5698, 159.7409, 
    161.9228, 164.1142, 166.3139, 168.5203, 170.7322, 172.9479, 175.166, 
    177.3849, 179.603, -178.1811, -175.9691, -173.7622, -171.5619, -169.3695, 
    -167.1861, -165.013, -162.8511, -160.7013, -158.5643, -156.4409, 
    -154.3314, -152.2363, -150.1559, -148.0902, -146.0393, -144.0032, 
    -141.9815, -139.9741, -137.9805, -136.0002, -134.0328, -132.0775, 
    -130.1339, -128.201, -126.2782, -124.3648, -122.4599, -120.5628, 
    -118.6726, -116.7887, -114.9103, -113.0367, -111.1671, -109.3009, 
    -107.4375, -105.5762, -103.7166, -101.858, -100, -98.14196, -96.28339, 
    -94.42377, -92.56254, -90.69913, -88.83294, -86.96335, -85.08969, 
    -83.21127, -81.32737, -79.43725, -77.54013, -75.63524, -73.72179, 
    -71.79903, -69.86616, -67.92245, -65.96722, -63.99977, -62.01952, 
    -60.02591, -58.01847, -55.99683, -53.96067, -51.90981, -49.84414, 
    -47.76369, -45.6686, -43.55913, -41.43565, -39.29869, -37.14887, 
    -34.98697, -32.81386, -30.63054, -28.43813, -26.23783, -24.03095, 
    -21.81886, -19.603, -17.38487, -15.16599, -12.94791, -10.73218, 
    -8.520334, -6.313863, -4.114222, -1.922801, 0.2590871, 2.430221, 
    4.589478, 6.735849, 8.868441, 10.98649, 13.08935, 15.17652, 17.24764, 
    19.30246, 21.34089, 23.36295, 25.3688, 27.35872, 29.33312, 31.29249, 
    33.23748, 35.16879, 37.08723, 38.99372, 40.88923, 42.77481, 44.65155, 
    46.52063, 48.38321, 50.24052, 52.09375, 53.94413, 55.79282, 57.64092, 
    59.48949, 61.33944, 63.19157, 65.04654, 66.90479, 68.76659, 70.632, 
    72.50081, 74.37267, 76.24699, 78.12305, 80,
  78.13536, 80, 81.86464, 83.72806, 85.5891, 87.44679, 89.30035, 91.14928, 
    92.99333, 94.83257, 96.66733, 98.49818, 100.326, 102.1516, 103.9763, 
    105.8014, 107.6281, 109.4578, 111.292, 113.1322, 114.9797, 116.8359, 
    118.7022, 120.5799, 122.4701, 124.3741, 126.2929, 128.2274, 130.1785, 
    132.1469, 134.1332, 136.1379, 138.1615, 140.2039, 142.2655, 144.346, 
    146.4452, 148.5627, 150.698, 152.8503, 155.0187, 157.2023, 159.3999, 
    161.6102, 163.8316, 166.0629, 168.3022, 170.5479, 172.7982, 175.0513, 
    177.3053, 179.5586, -178.1909, -175.9447, -173.7047, -171.4725, 
    -169.2495, -167.0372, -164.8369, -162.6499, -160.4769, -158.3191, 
    -156.1771, -154.0514, -151.9426, -149.8508, -147.7762, -145.7189, 
    -143.6786, -141.6552, -139.6482, -137.6572, -135.6817, -133.7208, 
    -131.774, -129.8405, -127.9193, -126.0097, -124.1107, -122.2215, 
    -120.3411, -118.4686, -116.6032, -114.7439, -112.8899, -111.0405, 
    -109.1949, -107.3523, -105.5122, -103.6738, -101.8366, -100, -98.16338, 
    -96.32618, -94.48782, -92.64767, -90.80513, -88.9595, -87.11008, 
    -85.25613, -83.39683, -81.53136, -79.65887, -77.77847, -75.88925, 
    -73.99029, -72.08069, -70.15955, -68.22598, -66.27918, -64.31835, 
    -62.34276, -60.35176, -58.34478, -56.32135, -54.2811, -52.22376, 
    -50.1492, -48.05743, -45.94858, -43.82292, -41.68089, -39.52306, 
    -37.35015, -35.16305, -32.96279, -30.75052, -28.52755, -26.29529, 
    -24.05528, -21.80914, -19.55857, -17.30535, -15.05127, -12.79817, 
    -10.54787, -8.302181, -6.062872, -3.831652, -1.610148, 0.6001045, 
    2.797682, 4.981283, 7.149745, 9.302042, 11.43731, 13.55482, 15.65402, 
    17.73451, 19.79605, 21.83854, 23.86206, 25.86681, 27.85314, 29.82153, 
    31.77261, 33.70711, 35.62587, 37.52985, 39.42011, 41.29779, 43.16409, 
    45.02031, 46.86781, 48.70796, 50.54219, 52.37193, 54.19862, 56.02365, 
    57.84837, 59.67405, 61.50182, 63.33267, 65.16743, 67.00667, 68.85072, 
    70.69965, 72.55321, 74.4109, 76.27194, 78.13536, 80,
  78.14803, 80, 81.85197, 83.70231, 85.54948, 87.39216, 89.22935, 91.06039, 
    92.88502, 94.70329, 96.51567, 98.3229, 100.126, 101.9262, 103.7249, 
    105.5236, 107.324, 109.1277, 110.9363, 112.7516, 114.5752, 116.4087, 
    118.2536, 120.1115, 121.9838, 123.8716, 125.7764, 127.6991, 129.6409, 
    131.6024, 133.5845, 135.5878, 137.6126, 139.6593, 141.7281, 143.8187, 
    145.931, 148.0645, 150.2187, 152.3927, 154.5856, 156.7962, 159.0231, 
    161.265, 163.52, 165.7865, 168.0625, 170.346, 172.635, 174.9274, 
    177.2209, 179.5134, -178.1972, -175.9129, -173.6359, -171.368, -169.1109, 
    -166.8664, -164.636, -162.421, -160.2226, -158.0418, -155.8794, 
    -153.7361, -151.6123, -149.5083, -147.4243, -145.3602, -143.3159, 
    -141.2909, -139.2848, -137.2971, -135.3271, -133.374, -131.4369, 
    -129.5149, -127.607, -125.7122, -123.8295, -121.9578, -120.0961, 
    -118.2432, -116.3983, -114.5602, -112.7281, -110.901, -109.078, 
    -107.2585, -105.4416, -103.6267, -101.813, -100, -98.18696, -96.37329, 
    -94.55836, -92.74148, -90.92196, -89.09904, -87.27194, -85.4398, 
    -83.60173, -81.75676, -79.90392, -78.04217, -76.17047, -74.28777, 
    -72.39301, -70.48514, -68.56314, -66.62604, -64.6729, -62.70287, 
    -60.71518, -58.70913, -56.68415, -54.63977, -52.57568, -50.49166, 
    -48.3877, -46.26392, -44.1206, -41.95821, -39.7774, -37.57899, -35.36399, 
    -33.13357, -30.88909, -28.63204, -26.36411, -24.08707, -21.80284, 
    -19.51342, -17.22089, -14.92738, -12.63505, -10.34604, -8.062498, 
    -5.786484, -3.520002, -1.264957, 0.9768662, 3.203821, 5.414408, 7.607293, 
    9.781315, 11.9355, 14.06904, 16.18133, 18.27194, 20.34065, 22.38737, 
    24.41223, 26.41549, 28.3976, 30.35915, 32.30086, 34.2236, 36.12836, 
    38.01624, 39.88847, 41.74636, 43.5913, 45.42479, 47.24838, 49.06367, 
    50.87231, 52.67598, 54.47635, 56.27509, 58.0738, 59.874, 61.6771, 
    63.48433, 65.29671, 67.11498, 68.93961, 70.77065, 72.60784, 74.45052, 
    76.29769, 78.14803, 80,
  78.16101, 80, 81.83899, 83.67581, 85.50845, 87.3352, 89.15477, 90.96635, 
    92.76962, 94.56475, 96.35233, 98.13334, 99.90905, 101.681, 103.4509, 
    105.2205, 106.9918, 108.7667, 110.5471, 112.335, 114.1323, 115.9407, 
    117.7621, 119.5982, 121.4505, 123.3206, 125.2098, 127.1194, 129.0506, 
    131.0044, 132.9816, 134.9829, 137.0089, 139.06, 141.1363, 143.2377, 
    145.3642, 147.5152, 149.6901, 151.888, 154.1078, 156.3482, 158.6077, 
    160.8846, 163.177, 165.4828, 167.7997, 170.1256, 172.4579, 174.7941, 
    177.1317, 179.4682, -178.199, -175.8722, -173.5538, -171.2461, -168.9512, 
    -166.6709, -164.4071, -162.1613, -159.9348, -157.7288, -155.5442, 
    -153.3817, -151.2418, -149.1248, -147.0309, -144.9598, -142.9114, 
    -140.8852, -138.8807, -136.8972, -134.9337, -132.9895, -131.0636, 
    -129.1547, -127.2618, -125.3837, -123.5192, -121.6671, -119.8261, 
    -117.995, -116.1728, -114.3581, -112.5501, -110.7476, -108.9497, 
    -107.1555, -105.3642, -103.575, -101.7872, -100, -98.21284, -96.42501, 
    -94.6358, -92.84448, -91.05029, -89.2524, -87.4499, -85.64185, -83.82723, 
    -82.00497, -80.17393, -78.33294, -76.4808, -74.61629, -72.7382, 
    -70.84531, -68.93645, -67.01045, -65.06626, -63.10284, -61.11929, 
    -59.11478, -57.0886, -55.04019, -52.96913, -50.87515, -48.75817, 
    -46.61829, -44.45579, -42.27119, -40.06519, -37.8387, -35.59288, 
    -33.32906, -31.04881, -28.75387, -26.44618, -24.12782, -21.80103, 
    -19.46817, -17.13168, -14.79406, -12.45785, -10.12558, -7.799734, 
    -5.482753, -3.176971, -0.8846001, 1.392291, 3.651803, 5.89222, 8.112026, 
    10.30991, 12.48479, 14.63579, 16.76225, 18.86374, 20.94002, 22.99109, 
    25.01711, 27.01844, 28.99563, 30.94939, 32.88058, 34.7902, 36.67941, 
    38.54948, 40.40179, 42.23787, 44.05928, 45.86774, 47.665, 49.4529, 
    51.23333, 53.00821, 54.7795, 56.54913, 58.31901, 60.09095, 61.86666, 
    63.64767, 65.43525, 67.23038, 69.03365, 70.84523, 72.6648, 74.49155, 
    76.32419, 78.16101, 80,
  78.17429, 80, 81.82571, 83.64857, 85.46597, 87.27575, 89.07627, 90.86657, 
    92.64633, 94.41584, 96.17593, 97.92784, 99.67321, 101.4139, 103.1519, 
    104.8895, 106.6288, 108.3721, 110.1216, 111.8795, 113.6479, 115.429, 
    117.2246, 119.0368, 120.8672, 122.7177, 124.5897, 126.4847, 128.4041, 
    130.349, 132.3205, 134.3194, 136.3463, 138.4017, 140.4859, 142.599, 
    144.7407, 146.9106, 149.1081, 151.3321, 153.5815, 155.8548, 158.1503, 
    160.4661, 162.7999, 165.1495, 167.5121, 169.8852, 172.2658, 174.651, 
    177.038, 179.4236, -178.195, -175.8207, -173.4563, -171.1044, -168.7673, 
    -166.4475, -164.1467, -161.867, -159.6097, -157.3762, -155.1674, 
    -152.9842, -150.8271, -148.6963, -146.5919, -144.5138, -142.4616, 
    -140.4347, -138.4325, -136.4541, -134.4985, -132.5647, -130.6514, 
    -128.7574, -126.8814, -125.022, -123.1778, -121.3474, -119.5294, 
    -117.7225, -115.9253, -114.1366, -112.355, -110.5796, -108.8091, 
    -107.0427, -105.2794, -103.5184, -101.7588, -100, -98.24117, -96.48161, 
    -94.72057, -92.95727, -91.19086, -89.42042, -87.64497, -85.86344, 
    -84.07469, -82.2775, -80.47058, -78.65262, -76.82223, -74.97803, 
    -73.11861, -71.24258, -69.34859, -67.43532, -65.50148, -63.54591, 
    -61.5675, -59.56529, -57.53842, -55.48619, -53.40807, -51.3037, 
    -49.17291, -47.01578, -44.83258, -42.62383, -40.3903, -38.13301, 
    -35.85325, -33.55254, -31.23265, -28.89563, -26.54368, -24.17927, 
    -21.80499, -19.4236, -17.03798, -14.65105, -12.26579, -9.885174, 
    -7.512117, -5.149462, -2.799928, -0.4660825, 1.849689, 4.145206, 
    6.418517, 8.66791, 10.89193, 13.08936, 15.25928, 17.40099, 19.51406, 
    21.5983, 23.65374, 25.68065, 27.67951, 29.65098, 31.5959, 33.51529, 
    35.41034, 37.28235, 39.13279, 40.96323, 42.77538, 44.57102, 46.35206, 
    48.1205, 49.8784, 51.62789, 53.37118, 55.11049, 56.84806, 58.5861, 
    60.32679, 62.07215, 63.82408, 65.58416, 67.35367, 69.13343, 70.92373, 
    72.72425, 74.53403, 76.35143, 78.17429, 80,
  78.18787, 80, 81.81213, 83.62057, 85.42197, 87.21355, 88.99336, 90.76028, 
    92.51405, 94.25517, 95.98476, 97.70447, 99.41631, 101.1225, 102.8256, 
    104.528, 106.2323, 107.9411, 109.6569, 111.3821, 113.1192, 114.8703, 
    116.6379, 118.4239, 120.2304, 122.0593, 123.9124, 125.7912, 127.6975, 
    129.6324, 131.5972, 133.5928, 135.6203, 137.68, 139.7725, 141.8978, 
    144.0558, 146.2461, 148.4681, 150.7206, 153.0024, 155.3119, 157.6472, 
    160.006, 162.3858, 164.7841, 167.1976, 169.6234, 172.058, 174.498, 
    176.9401, 179.3806, -178.1838, -175.7565, -173.3408, -170.9397, -168.556, 
    -166.1922, -163.8508, -161.5338, -159.2428, -156.9793, -154.7444, 
    -152.539, -150.3635, -148.2182, -146.1032, -144.018, -141.9624, 
    -139.9355, -137.9365, -135.9645, -134.0182, -132.0963, -130.1975, 
    -128.3204, -126.4633, -124.6248, -122.8031, -120.9969, -119.2044, 
    -117.4241, -115.6545, -113.8942, -112.1418, -110.396, -108.6556, 
    -106.9196, -105.1869, -103.4566, -101.7279, -100, -98.27209, -96.5434, 
    -94.81313, -93.08044, -91.34441, -89.60404, -87.85824, -86.10582, 
    -84.3455, -82.57591, -80.79562, -79.00312, -77.19685, -75.37524, 
    -73.5367, -71.67963, -69.80247, -67.90369, -65.98183, -64.03552, 
    -62.06347, -60.06452, -58.03764, -55.98197, -53.89684, -51.78176, 
    -49.63649, -47.46101, -45.25557, -43.02069, -40.75721, -38.46622, 
    -36.14916, -33.80776, -31.44404, -29.06031, -26.65917, -24.24345, 
    -21.81618, -19.38061, -16.94007, -14.49803, -12.05796, -9.623345, 
    -7.197607, -4.784056, -2.385854, -0.005973984, 2.352843, 4.688106, 
    6.997604, 9.279421, 11.53194, 13.75386, 15.94418, 18.10219, 20.2275, 
    22.31997, 24.37972, 26.40714, 28.40284, 30.36764, 32.30254, 34.20876, 
    36.08764, 37.94069, 39.76958, 41.57609, 43.36211, 45.12965, 46.88084, 
    48.61789, 50.34311, 52.05888, 53.76767, 55.47199, 57.1744, 58.87746, 
    60.5837, 62.29553, 64.01524, 65.74483, 67.48595, 69.23972, 71.00664, 
    72.78645, 74.57803, 76.37943, 78.18787, 80,
  78.20172, 80, 81.79828, 83.59179, 85.37626, 87.14825, 88.9054, 90.6465, 
    92.37144, 94.08105, 95.77684, 97.46095, 99.13584, 100.8043, 102.469, 
    104.1331, 105.7994, 107.4707, 109.1499, 110.8397, 112.5427, 114.2616, 
    115.9986, 117.7562, 119.5366, 121.3419, 123.1741, 125.0351, 126.9266, 
    128.8501, 130.8071, 132.7988, 134.8262, 136.89, 138.9909, 141.129, 
    143.3043, 145.5165, 147.7649, 150.0484, 152.3656, 154.7148, 157.0939, 
    159.5003, 161.9313, 164.3836, 166.8538, 169.3384, 171.8333, 174.3346, 
    176.8383, 179.3402, -178.1636, -175.6773, -173.2044, -170.7486, 
    -168.3131, -165.9009, -163.5147, -161.1568, -158.829, -156.5331, 
    -154.2701, -152.0409, -149.846, -147.6857, -145.5597, -143.4678, 
    -141.4093, -139.3833, -137.3888, -135.4246, -133.4892, -131.5811, 
    -129.6989, -127.8407, -126.0049, -124.1896, -122.3931, -120.6135, 
    -118.8491, -117.0981, -115.3588, -113.6297, -111.9091, -110.1958, 
    -108.4882, -106.7854, -105.0861, -103.3893, -101.6942, -100, -98.30576, 
    -96.61069, -94.91395, -93.21465, -91.51177, -89.80424, -88.09085, 
    -86.3703, -84.64115, -82.90189, -81.15089, -79.38648, -77.6069, 
    -75.81038, -73.9951, -72.15927, -70.3011, -68.41885, -66.51083, 
    -64.57544, -62.61118, -60.61667, -58.59068, -56.53217, -54.44026, 
    -52.31433, -50.15399, -47.95913, -45.72995, -43.46695, -41.17097, 
    -38.84324, -36.4853, -34.09909, -31.68693, -29.25144, -26.79562, 
    -24.32274, -21.83636, -19.34025, -16.83833, -14.33465, -11.8333, 
    -9.338361, -6.853831, -4.383572, -1.931257, 0.4996836, 2.906103, 
    5.285168, 7.63439, 9.951635, 12.23514, 14.4835, 16.69569, 18.87101, 
    21.00911, 23.10996, 25.1738, 27.20118, 29.19287, 31.14988, 33.07342, 
    34.9649, 36.82587, 38.65808, 40.46339, 42.24379, 44.00139, 45.73844, 
    47.45726, 49.1603, 50.8501, 52.5293, 54.20063, 55.8669, 57.53096, 
    59.19575, 60.86416, 62.53905, 64.22316, 65.91895, 67.62856, 69.3535, 
    71.0946, 72.85175, 74.62374, 76.40821, 78.20172, 80,
  78.21587, 80, 81.78413, 83.56214, 85.32861, 87.07931, 88.8115, 90.52396, 
    92.21687, 93.89146, 95.54986, 97.19472, 98.82907, 100.4562, 102.0793, 
    103.7017, 105.3268, 106.9577, 108.5974, 110.2491, 111.9154, 113.5993, 
    115.3034, 117.0302, 118.7822, 120.5617, 122.371, 124.2122, 126.0871, 
    127.9978, 129.9456, 131.9323, 133.9588, 136.0264, 138.1355, 140.2869, 
    142.4804, 144.7158, 146.9926, 149.3097, 151.6655, 154.0582, 156.4855, 
    158.9445, 161.4321, 163.9445, 166.478, 169.0282, 171.5906, 174.1605, 
    176.7332, 179.3038, -178.1324, -175.58, -173.0435, -170.5269, -168.0341, 
    -165.5684, -163.1329, -160.7303, -158.3626, -156.0315, -153.7384, 
    -151.484, -149.2689, -147.0931, -144.9564, -142.8582, -140.7976, 
    -138.7737, -136.7851, -134.8303, -132.9078, -131.0157, -129.1523, 
    -127.3155, -125.5034, -123.7141, -121.9453, -120.1952, -118.4617, 
    -116.7428, -115.0368, -113.3417, -111.656, -109.9779, -108.3062, 
    -106.6394, -104.9764, -103.3162, -101.6577, -100, -98.34235, -96.68383, 
    -95.02357, -93.36057, -91.6938, -90.02206, -88.34402, -86.65827, 
    -84.96321, -83.25716, -81.53833, -79.80482, -78.0547, -76.28595, 
    -74.49656, -72.68449, -70.84772, -68.98427, -67.0922, -65.16966, 
    -63.2149, -61.2263, -59.20237, -57.14185, -55.04364, -52.90691, 
    -50.73111, -48.51598, -46.26162, -43.96848, -41.63742, -39.26971, 
    -36.86705, -34.43161, -31.96595, -29.4731, -26.95651, -24.41995, 
    -21.86757, -19.30377, -16.73317, -14.1605, -11.59058, -9.028193, 
    -6.478014, -3.944551, -1.432066, 1.055483, 3.514496, 5.94176, 8.33449, 
    10.69033, 13.00738, 15.28416, 17.51963, 19.71314, 21.86445, 23.97365, 
    26.04117, 28.06774, 30.05435, 32.00224, 33.91286, 35.78784, 37.629, 
    39.4383, 41.21784, 42.96984, 44.69664, 46.4007, 48.08458, 49.75094, 
    51.40256, 53.04231, 54.67318, 56.29825, 57.92072, 59.54384, 61.17093, 
    62.80528, 64.45014, 66.10854, 67.78313, 69.47604, 71.1885, 72.92069, 
    74.67139, 76.43786, 78.21587, 80,
  78.23033, 80, 81.76967, 83.53151, 85.27869, 87.00607, 88.71057, 90.39113, 
    92.04833, 93.68408, 95.30116, 96.90292, 98.493, 100.0752, 101.6532, 
    103.2308, 104.8115, 106.3989, 107.9963, 109.6069, 111.2339, 112.8802, 
    114.5487, 116.2422, 117.9634, 119.7148, 121.4989, 123.3181, 125.1746, 
    127.0705, 129.0077, 130.9878, 133.0126, 135.0831, 137.2004, 139.3651, 
    141.5775, 143.8376, 146.1447, 148.4979, 150.8956, 153.3359, 155.8161, 
    158.3332, 160.8835, 163.4629, 166.0669, 168.6904, 171.3284, 173.9751, 
    176.6251, 179.2727, -178.0878, -175.4616, -172.854, -170.2699, -167.7135, 
    -165.1888, -162.6993, -160.2478, -157.8368, -155.468, -153.1428, 
    -150.8619, -148.6258, -146.4344, -144.2872, -142.1834, -140.1221, 
    -138.1017, -136.1208, -134.1776, -132.2701, -130.3964, -128.5543, 
    -126.7416, -124.9561, -123.1954, -121.4574, -119.7396, -118.0401, 
    -116.3564, -114.6867, -113.0288, -111.381, -109.7414, -108.1086, 
    -106.481, -104.8575, -103.2368, -101.618, -100, -98.38205, -96.76321, 
    -95.14252, -93.51897, -91.89143, -90.25858, -88.61904, -86.97119, 
    -85.31333, -83.64357, -81.95995, -80.26035, -78.54265, -76.8046, 
    -75.04395, -73.25841, -71.44572, -69.60361, -67.7299, -65.82246, 
    -63.87922, -61.89831, -59.87794, -57.81656, -55.71282, -53.56562, 
    -51.37419, -49.13808, -46.85723, -44.53199, -42.1632, -39.75216, 
    -37.3007, -34.81119, -32.28652, -29.73013, -27.14596, -24.53839, 
    -21.91224, -19.27268, -16.62511, -13.97512, -11.32836, -8.690451, 
    -6.066887, -3.462926, -0.8835167, 1.666781, 4.183854, 6.664079, 9.104353, 
    11.50211, 13.85531, 16.16244, 18.4225, 20.63493, 22.79964, 24.91693, 
    26.98744, 29.01216, 30.99234, 32.92951, 34.82539, 36.68188, 38.50108, 
    40.28522, 42.03663, 43.7578, 45.45129, 47.11979, 48.76609, 50.39305, 
    52.00368, 53.60108, 55.18848, 56.76923, 58.34682, 59.92484, 61.507, 
    63.09708, 64.69884, 66.31592, 67.95167, 69.60887, 71.28943, 72.99393, 
    74.72131, 76.46849, 78.23033, 80,
  78.24512, 80, 81.75488, 83.49973, 85.22602, 86.92762, 88.60122, 90.24609, 
    91.8635, 93.45621, 95.02782, 96.58247, 98.12443, 99.65804, 101.1875, 
    102.717, 104.2503, 105.7912, 107.3434, 108.9102, 110.495, 112.101, 
    113.7312, 115.3888, 117.0765, 118.7973, 120.5537, 122.3486, 124.1843, 
    126.0633, 127.9878, 129.9599, 131.9813, 134.0538, 136.1786, 138.3566, 
    140.5884, 142.8742, 145.2135, 147.6055, 150.0486, 152.5407, 155.079, 
    157.6601, 160.28, 162.9339, 165.6166, 168.3223, 171.0449, 173.7779, 
    176.5148, 179.2487, -178.0267, -175.318, -172.6311, -169.9718, -167.345, 
    -164.7553, -162.2065, -159.7019, -157.244, -154.8349, -152.4757, 
    -150.1672, -147.9097, -145.7027, -143.5458, -141.4376, -139.377, 
    -137.362, -135.391, -133.4617, -131.5719, -129.7193, -127.9014, 
    -126.1157, -124.3598, -122.631, -120.9267, -119.2446, -117.5822, 
    -115.937, -114.3068, -112.6894, -111.0828, -109.485, -107.8944, 
    -106.3094, -104.7286, -103.1508, -101.5749, -100, -98.42507, -96.84921, 
    -95.27142, -93.69064, -92.10562, -90.515, -88.91724, -87.3106, -85.6932, 
    -84.063, -82.41782, -80.75536, -79.07326, -77.36905, -75.64023, 
    -73.88426, -72.0986, -70.28072, -68.42811, -66.53834, -64.60904, 
    -62.63797, -60.62305, -58.56236, -56.45423, -54.29725, -52.09034, 
    -49.83279, -47.52431, -45.16513, -42.75595, -40.2981, -37.79351, 
    -35.24474, -32.65501, -30.02821, -27.36884, -24.682, -21.97329, 
    -19.24875, -16.51477, -13.77793, -11.04489, -8.322294, -5.616578, 
    -2.933898, -0.2800027, 2.339852, 4.920978, 7.459304, 9.951404, 12.3945, 
    14.78646, 17.12579, 19.41156, 21.64339, 23.82142, 25.94619, 28.01866, 
    30.04014, 32.0122, 33.93671, 35.8157, 37.65143, 39.44627, 41.20274, 
    42.92348, 44.61122, 46.26876, 47.89902, 49.50501, 51.08982, 52.65664, 
    54.2088, 55.74973, 57.28304, 58.81248, 60.34196, 61.87557, 63.41753, 
    64.97218, 66.54379, 68.1365, 69.75391, 71.39878, 73.07238, 74.77398, 
    76.50027, 78.24512, 80,
  78.26032, 80, 81.73968, 83.46656, 85.16999, 86.84283, 88.48172, 90.08657, 
    91.65968, 93.20483, 94.72665, 96.23007, 97.72008, 99.20152, 100.6791, 
    102.1572, 103.64, 105.1315, 106.6355, 108.1557, 109.6955, 111.2584, 
    112.8476, 114.4664, 116.1179, 117.8052, 119.5313, 121.299, 123.1113, 
    124.9709, 126.8804, 128.8423, 130.8587, 132.9316, 135.0629, 137.2537, 
    139.5051, 141.8174, 144.1906, 146.6239, 149.1158, 151.6642, 154.2662, 
    156.9179, 159.6149, 162.3518, 165.1225, 167.9203, 170.7381, 173.5683, 
    176.4029, 179.2341, -177.9458, -175.1445, -172.369, -169.6259, -166.9211, 
    -164.2597, -161.646, -159.0837, -156.5755, -154.1234, -151.7286, 
    -149.3917, -147.1126, -144.8907, -142.7251, -140.6142, -138.5562, 
    -136.5491, -134.5905, -132.678, -130.8089, -128.9805, -127.19, -125.4347, 
    -123.7116, -122.018, -120.351, -118.7078, -117.0859, -115.4826, 
    -113.8954, -112.3219, -110.76, -109.2075, -107.6626, -106.1236, 
    -104.5891, -103.0577, -101.5284, -100, -98.47163, -96.94227, -95.41091, 
    -93.87639, -92.33743, -90.79253, -89.24003, -87.67806, -86.10458, 
    -84.51737, -82.91405, -81.29215, -79.64904, -77.98205, -76.28841, 
    -74.56534, -72.80999, -71.01953, -69.19114, -67.32204, -65.4095, 
    -63.45091, -61.44378, -59.3858, -57.27489, -55.10925, -52.88742, 
    -50.60833, -48.2714, -45.87659, -43.42447, -40.91627, -38.35398, 
    -35.74035, -33.07893, -30.37409, -27.63098, -24.8555, -22.05418, 
    -19.23414, -16.4029, -13.56827, -10.73813, -7.920329, -5.122468, 
    -2.351758, 0.3851079, 3.082079, 5.733824, 8.335783, 10.88421, 13.37614, 
    15.80941, 18.18258, 20.49492, 22.74629, 24.93713, 27.06837, 29.14133, 
    31.15774, 33.11956, 35.02906, 36.88866, 38.70098, 40.46874, 42.1948, 
    43.88208, 45.53357, 47.15237, 48.7416, 50.30449, 51.84432, 53.3645, 
    54.86853, 56.36004, 57.84285, 59.32092, 60.79848, 62.27992, 63.76993, 
    65.27335, 66.79517, 68.34032, 69.91343, 71.51828, 73.15717, 74.83001, 
    76.53344, 78.26032, 80,
  78.27597, 80, 81.72403, 83.43168, 85.10979, 86.75024, 88.34995, 89.90994, 
    91.43383, 92.92671, 94.39429, 95.84238, 97.27663, 98.7024, 100.1247, 
    101.5483, 102.9777, 104.4168, 105.8699, 107.3406, 108.8326, 110.3495, 
    111.8947, 113.4718, 115.0841, 116.7348, 118.4274, 120.165, 121.9508, 
    123.7881, 125.6797, 127.6287, 129.6376, 131.7091, 133.8452, 136.0479, 
    138.3184, 140.6578, 143.0661, 145.5431, 148.0873, 150.6968, 153.3683, 
    156.0978, 158.8803, 161.7097, 164.579, 167.4805, 170.4056, 173.3453, 
    176.2904, 179.2314, -177.8409, -174.9354, -172.0607, -169.2242, 
    -166.4328, -163.6925, -161.008, -158.3833, -155.8212, -153.3237, 
    -150.8919, -148.5261, -146.2258, -143.9902, -141.8176, -139.7061, 
    -137.6534, -135.657, -133.714, -131.8216, -129.9766, -128.1759, 
    -126.4165, -124.6951, -123.0085, -121.3537, -119.7275, -118.127, 
    -116.5492, -114.9914, -113.4508, -111.9248, -110.4112, -108.9076, 
    -107.4121, -105.9229, -104.4383, -102.9571, -101.4781, -100, -98.52193, 
    -97.04285, -95.56166, -94.07714, -92.58792, -91.09242, -89.58884, 
    -88.07519, -86.54925, -85.00863, -83.45079, -81.87302, -80.27251, 
    -78.64635, -76.99152, -75.30495, -73.58351, -71.82406, -70.02342, 
    -68.17844, -66.28598, -64.343, -62.34657, -60.29389, -58.1824, -56.0098, 
    -53.77415, -51.47392, -49.10811, -46.67632, -44.17883, -41.61675, 
    -38.99202, -36.30753, -33.56717, -30.77581, -27.93934, -25.06456, 
    -22.15913, -19.23145, -16.29042, -13.34533, -10.40558, -7.48047, 
    -4.57901, -1.709686, 1.119708, 3.902194, 6.631727, 9.303235, 11.91266, 
    14.45691, 16.93385, 19.34223, 21.68158, 23.95215, 26.1548, 28.29094, 
    30.36238, 32.37133, 34.32027, 36.21192, 38.04916, 39.83503, 41.57264, 
    43.2652, 44.91595, 46.52819, 48.10526, 49.65053, 51.16743, 52.65944, 
    54.13012, 55.58316, 57.02235, 58.45166, 59.87526, 61.2976, 62.72338, 
    64.15762, 65.60571, 67.07329, 68.56617, 70.09006, 71.65005, 73.24976, 
    74.89021, 76.56832, 78.27597, 80,
  78.29219, 80, 81.70781, 83.39465, 85.04436, 86.64801, 88.20341, 89.71317, 
    91.18262, 92.61837, 94.02728, 95.41602, 96.79088, 98.15762, 99.52161, 
    100.8878, 102.2607, 103.6447, 105.0439, 106.4623, 107.9035, 109.3715, 
    110.8697, 112.4019, 113.9716, 115.5824, 117.238, 118.942, 120.6979, 
    122.5093, 124.3797, 126.3125, 128.3109, 130.3781, 132.5169, 134.7297, 
    137.0185, 139.3847, 141.8292, 144.3519, 146.9518, 149.627, 152.3743, 
    155.1894, 158.0668, 160.9995, 163.9795, 166.9978, 170.0442, 173.1082, 
    176.1785, 179.2439, -177.7067, -174.6839, -171.6977, -168.757, -165.8697, 
    -163.0425, -160.2808, -157.5887, -154.9694, -152.4244, -149.9548, 
    -147.5602, -145.2399, -142.9922, -140.8151, -138.7059, -136.6618, 
    -134.6796, -132.756, -130.8875, -129.0706, -127.3017, -125.5773, 
    -123.8937, -122.2476, -120.6354, -119.0539, -117.4998, -115.9699, 
    -114.4613, -112.9711, -111.4964, -110.0348, -108.584, -107.1417, 
    -105.7062, -104.2756, -102.8485, -101.4237, -100, -98.57626, -97.15145, 
    -95.7244, -94.29382, -92.85825, -91.416, -89.96516, -88.50359, -87.02895, 
    -85.53867, -84.03005, -82.5002, -80.94608, -79.36458, -77.75243, 
    -76.10629, -74.42274, -72.69827, -70.92937, -69.11246, -67.24397, 
    -65.32037, -63.33818, -61.29409, -59.18492, -57.00777, -54.7601, 
    -52.43978, -50.04523, -47.57556, -45.03064, -42.41125, -39.71924, 
    -36.95754, -34.13033, -31.24302, -28.3023, -25.31605, -22.29326, 
    -19.24385, -16.17845, -13.10815, -10.04421, -6.997763, -3.979512, 
    -0.9994779, 1.933225, 4.810559, 7.625686, 10.37301, 13.0482, 15.64812, 
    18.1708, 20.61527, 22.98152, 25.27031, 27.48308, 29.62185, 31.68907, 
    33.68753, 35.62032, 37.49071, 39.3021, 41.058, 42.76196, 44.41757, 
    46.02843, 47.59814, 49.13031, 50.62854, 52.09646, 53.53773, 54.95607, 
    56.35528, 57.7393, 59.11223, 60.47839, 61.84238, 63.20913, 64.58398, 
    65.97272, 67.38163, 68.81738, 70.28683, 71.79659, 73.35199, 74.95564, 
    76.60535, 78.29219, 80,
  78.3091, 80, 81.6909, 83.35486, 84.9723, 86.53391, 88.03915, 89.49286, 
    90.9025, 92.27628, 93.62225, 94.94785, 96.25987, 97.56445, 98.86715, 
    100.173, 101.4868, 102.8129, 104.1555, 105.5186, 106.9062, 108.322, 
    109.77, 111.2539, 112.7775, 114.3447, 115.9596, 117.6259, 119.3478, 
    121.1292, 122.9743, 124.8869, 126.871, 128.9305, 131.0688, 133.2891, 
    135.5943, 137.9865, 140.4673, 143.0373, 145.6959, 148.4416, 151.2713, 
    154.1805, 157.163, 160.2112, 163.3158, 166.4662, 169.6503, 172.8555, 
    176.0684, 179.2753, -177.5372, -174.3816, -171.2699, -168.2127, 
    -165.2189, -162.2963, -159.4508, -156.6866, -154.0069, -151.4129, 
    -148.9052, -146.4828, -144.1443, -141.8873, -139.7089, -137.6059, 
    -135.5744, -133.6108, -131.7111, -129.871, -128.0867, -126.354, -124.669, 
    -123.0276, -121.4261, -119.8608, -118.328, -116.8243, -115.3462, 
    -113.8907, -112.4547, -111.0352, -109.6296, -108.2354, -106.8504, 
    -105.4726, -104.1001, -102.7314, -101.3651, -100, -98.63488, -97.26859, 
    -95.89989, -94.5274, -93.14956, -91.76457, -90.37041, -88.96484, 
    -87.54535, -86.10928, -84.65376, -83.17572, -81.67198, -80.13919, 
    -78.57386, -76.97238, -75.33102, -73.64597, -71.91328, -70.12895, 
    -68.28894, -66.38917, -64.42557, -62.39415, -60.29107, -58.11269, 
    -55.85569, -53.51719, -51.09485, -48.58708, -45.99314, -43.31335, 
    -40.54923, -37.70367, -34.78104, -31.78732, -28.73006, -25.61838, 
    -22.46284, -19.27526, -16.06837, -12.85554, -9.650334, -6.466154, 
    -3.315815, -0.2112067, 2.836993, 5.819531, 8.728698, 11.55839, 14.30408, 
    16.96273, 19.53267, 22.01346, 24.40571, 26.71089, 28.93123, 31.06951, 
    33.12895, 35.1131, 37.02573, 38.87076, 40.6522, 42.37407, 44.04042, 
    45.65525, 47.22252, 48.74615, 50.23002, 51.67796, 53.0938, 54.48135, 
    55.84447, 57.18707, 58.51317, 59.82696, 61.13285, 62.43555, 63.74013, 
    65.05215, 66.37775, 67.72372, 69.0975, 70.50714, 71.96085, 73.46609, 
    75.0277, 76.64514, 78.3091, 80,
  78.32689, 80, 81.67311, 83.31152, 84.89183, 86.40523, 87.85381, 89.24541, 
    90.58985, 91.89702, 93.17602, 94.43497, 95.68105, 96.92059, 98.15928, 
    99.40227, 100.6543, 101.9198, 103.203, 104.5081, 105.8389, 107.1994, 
    108.5936, 110.0256, 111.4993, 113.0189, 114.5887, 116.2129, 117.8961, 
    119.6428, 121.4576, 123.3452, 125.3103, 127.3574, 129.491, 131.7152, 
    134.0339, 136.4502, 138.9666, 141.5845, 144.3044, 147.1251, 150.0439, 
    153.0561, 156.1553, 159.3328, 162.5779, 165.8782, 169.2194, 172.586, 
    175.9619, 179.3305, -177.3244, -174.0181, -170.765, -167.5772, -164.4655, 
    -161.4383, -158.5021, -155.6613, -152.9185, -150.2748, -147.7296, 
    -145.2815, -142.9279, -140.6654, -138.4902, -136.398, -134.3843, 
    -132.4445, -130.5738, -128.7675, -127.0209, -125.3294, -123.6886, 
    -122.0942, -120.5419, -119.0277, -117.5479, -116.0986, -114.6765, 
    -113.278, -111.9, -110.5397, -109.194, -107.8606, -106.537, -105.2211, 
    -103.9111, -102.6052, -101.3019, -100, -98.69805, -97.39481, -96.08892, 
    -94.77888, -93.463, -92.1394, -90.80597, -89.46034, -88.09995, -86.72202, 
    -85.32355, -83.90137, -82.45212, -80.97227, -79.45813, -77.90584, 
    -76.31138, -74.67058, -72.9791, -71.2325, -69.42619, -67.55549, 
    -65.61567, -63.60201, -61.50983, -59.33461, -57.07211, -54.71846, 
    -52.27035, -49.72524, -47.08151, -44.33875, -41.49794, -38.56171, 
    -35.5345, -32.42279, -29.23505, -25.98185, -22.67564, -19.33053, 
    -15.96192, -12.58602, -9.219361, -5.878171, -2.577911, 0.6672379, 
    3.844726, 6.943903, 9.956149, 12.87491, 15.69559, 18.41547, 21.03344, 
    23.54982, 25.96611, 28.28477, 30.50901, 32.6426, 34.6897, 36.65476, 
    38.54237, 40.35719, 42.10388, 43.78708, 45.41133, 46.98109, 48.5007, 
    49.97441, 51.40635, 52.8006, 54.16114, 55.49195, 56.79696, 58.08018, 
    59.3457, 60.59773, 61.84072, 63.07941, 64.31895, 65.56503, 66.82398, 
    68.10298, 69.41015, 70.75459, 72.14619, 73.59477, 75.10817, 76.68848, 
    78.32689, 80,
  78.34581, 80, 81.65419, 83.26354, 84.80071, 86.25874, 87.64371, 88.96706, 
    90.24115, 91.47741, 92.68584, 93.87503, 95.05238, 96.22433, 97.39655, 
    98.5742, 99.76199, 100.9643, 102.1855, 103.4295, 104.7005, 106.0024, 
    107.3394, 108.7155, 110.1352, 111.6027, 113.1226, 114.6997, 116.339, 
    118.0454, 119.8242, 121.681, 123.6211, 125.6501, 127.7735, 129.9966, 
    132.3244, 134.7614, 137.3113, 139.9769, 142.7596, 145.6592, 148.6737, 
    151.7985, 155.0269, 158.3493, 161.7534, 165.2245, 168.7456, 172.2978, 
    175.8613, 179.4158, -177.0587, -173.5807, -170.1674, -166.8335, -163.591, 
    -160.4496, -157.4159, -154.4944, -151.687, -148.9939, -146.4136, 
    -143.9431, -141.5788, -139.316, -137.1497, -135.0745, -133.0848, 
    -131.175, -129.3395, -127.5728, -125.8697, -124.225, -122.6338, 
    -121.0913, -119.593, -118.1346, -116.7121, -115.3216, -113.9593, 
    -112.6219, -111.306, -110.0087, -108.727, -107.4583, -106.2003, 
    -104.9508, -103.7077, -102.4693, -101.2339, -100, -98.7661, -97.53071, 
    -96.2923, -95.04922, -93.79967, -92.54167, -91.27303, -89.99135, 
    -88.69399, -87.37813, -86.0407, -84.67844, -83.2879, -81.86538, 
    -80.40702, -78.90874, -77.36623, -75.77499, -74.13028, -72.42718, 
    -70.66054, -68.82504, -66.91522, -64.92551, -62.85027, -60.68396, 
    -58.42118, -56.05685, -53.58643, -51.00607, -48.31296, -45.50559, 
    -42.58406, -39.55042, -36.40897, -33.16654, -29.83258, -26.41927, 
    -22.94133, -19.41575, -15.86128, -12.29778, -8.745563, -5.224511, 
    -1.753403, 1.650725, 4.973094, 8.201474, 11.32632, 14.34075, 17.24039, 
    20.02309, 22.68869, 25.23861, 27.6756, 30.00341, 32.22652, 34.34992, 
    36.37893, 38.31903, 40.17577, 41.95464, 43.66105, 45.30026, 46.87739, 
    48.39734, 49.86484, 51.28447, 52.66064, 53.9976, 55.29953, 56.57048, 
    57.81451, 59.03565, 60.238, 61.4258, 62.60345, 63.77568, 64.94762, 
    66.12497, 67.31416, 68.52259, 69.75885, 71.03294, 72.35629, 73.74126, 
    75.19929, 76.73646, 78.34581, 80,
  78.36622, 80, 81.63378, 83.20947, 84.69615, 86.09082, 87.40499, 88.65418, 
    89.8532, 91.01477, 92.14952, 93.2663, 94.37255, 95.47466, 96.57824, 
    97.68833, 98.80956, 99.94629, 101.1027, 102.2829, 103.4908, 104.7307, 
    106.0066, 107.3229, 108.684, 110.0946, 111.5595, 113.0839, 114.6732, 
    116.333, 118.0692, 119.8881, 121.7962, 123.7999, 125.9061, 128.1213, 
    130.4522, 132.9047, 135.4844, 138.1955, 141.0412, 144.0228, 147.1391, 
    150.3863, 153.7575, 157.2423, 160.8268, 164.4934, 168.2217, 171.9885, 
    175.7692, 179.5387, -176.7278, -173.0533, -169.4584, -165.9604, 
    -162.5735, -159.3079, -156.1706, -153.1653, -150.2931, -147.5527, 
    -144.9411, -142.4536, -140.0849, -137.8288, -135.6787, -133.6279, 
    -131.6696, -129.7971, -128.0039, -126.2838, -124.6306, -123.0388, 
    -121.5028, -120.0177, -118.5785, -117.1806, -115.82, -114.4924, 
    -113.1941, -111.9217, -110.6717, -109.4413, -108.2274, -107.0276, 
    -105.8394, -104.6607, -103.4892, -102.3232, -101.1607, -100, -98.83929, 
    -97.67682, -96.51079, -95.33934, -94.16056, -92.97237, -91.77257, 
    -90.55874, -89.32827, -88.07835, -86.8059, -85.50764, -84.18005, 
    -82.81935, -81.42154, -79.98232, -78.49715, -76.96121, -75.36938, 
    -73.71623, -71.99606, -70.20287, -68.33037, -66.37206, -64.32127, 
    -62.17119, -59.91508, -57.54639, -55.05895, -52.44727, -49.70689, 
    -46.8347, -43.82944, -40.69212, -37.42652, -34.03956, -30.54162, 
    -26.94667, -23.27216, -19.53867, -15.76923, -11.98851, -8.221694, 
    -4.49344, -0.8267874, 2.757682, 6.242513, 9.613737, 12.86095, 15.97722, 
    18.95875, 21.80448, 24.51564, 27.09528, 29.54781, 31.87867, 34.09394, 
    36.20011, 38.20385, 40.11188, 41.9308, 43.66705, 45.32682, 46.91607, 
    48.44046, 49.90539, 51.31597, 52.67708, 53.99338, 55.26931, 56.50918, 
    57.71715, 58.89731, 60.05371, 61.19044, 62.31167, 63.42176, 64.52534, 
    65.62745, 66.7337, 67.85048, 68.98523, 70.1468, 71.34582, 72.59501, 
    73.90918, 75.30385, 76.79053, 78.36622, 80,
  78.38859, 80, 81.61141, 83.14738, 84.57478, 85.89749, 87.13382, 88.30347, 
    89.42335, 90.5071, 91.56566, 92.60787, 93.64105, 94.67144, 95.70446, 
    96.74499, 97.7975, 98.86626, 99.95534, 101.0688, 102.2106, 103.3849, 
    104.5959, 105.8481, 107.1459, 108.4944, 109.8986, 111.3641, 112.8967, 
    114.5027, 116.1886, 117.9616, 119.829, 121.7988, 123.8788, 126.0776, 
    128.4032, 130.8638, 133.4669, 136.2193, 139.1262, 142.1909, 145.4141, 
    148.7933, 152.3219, 155.9889, 159.7785, 163.67, 167.6384, 171.6552, 
    175.6894, 179.7092, -176.3163, -172.4157, -168.6141, -164.9323, 
    -161.3861, -157.9866, -154.7404, -151.6502, -148.7151, -145.9319, 
    -143.2953, -140.7985, -138.434, -136.1936, -134.069, -132.0518, 
    -130.1338, -128.3071, -126.5643, -124.8983, -123.3022, -121.7699, 
    -120.2954, -118.8732, -117.4984, -116.1659, -114.8716, -113.6112, 
    -112.3809, -111.1773, -109.997, -108.8371, -107.6949, -106.5678, 
    -105.4536, -104.35, -103.2549, -102.1663, -101.0821, -100, -98.91795, 
    -97.83369, -96.7451, -95.65005, -94.54645, -93.43221, -92.30513, 
    -91.1629, -90.00301, -88.82274, -87.61908, -86.38881, -85.1284, 
    -83.83405, -82.50165, -81.12675, -79.70462, -78.23013, -76.6978, 
    -75.10175, -73.43567, -71.69288, -69.86624, -67.94824, -65.931, 
    -63.80635, -61.56596, -59.20146, -56.70471, -54.06809, -51.2849, 
    -48.34983, -45.25956, -42.01337, -38.6139, -35.06771, -31.38589, 
    -27.58433, -23.68373, -19.7092, -15.68938, -11.65521, -7.638435, 
    -3.669986, 0.221544, 4.011128, 7.678132, 11.20674, 14.58592, 17.80915, 
    20.87385, 23.78072, 26.53309, 29.13624, 31.59684, 33.92245, 36.12115, 
    38.20124, 40.17097, 42.03843, 43.8114, 45.49734, 47.10329, 48.63589, 
    50.10138, 51.50561, 52.85408, 54.15195, 55.40409, 56.61512, 57.78942, 
    58.93124, 60.04467, 61.13374, 62.2025, 63.25502, 64.29554, 65.32856, 
    66.35895, 67.39213, 68.43434, 69.4929, 70.57665, 71.69653, 72.86618, 
    74.10251, 75.42522, 76.85262, 78.38859, 80,
  78.41363, 80, 81.58637, 83.07472, 84.43271, 85.67469, 86.82671, 87.91225, 
    88.94976, 89.95331, 90.93377, 91.89977, 92.85836, 93.81548, 94.7763, 
    95.74548, 96.72731, 97.72587, 98.74512, 99.78901, 100.8615, 101.9667, 
    103.1088, 104.2924, 105.5221, 106.8029, 108.1404, 109.5403, 111.0089, 
    112.553, 114.1799, 115.8976, 117.7144, 119.6396, 121.6827, 123.8538, 
    126.1632, 128.6215, 131.2389, 134.025, 136.9881, 140.1346, 143.468, 
    146.9879, 150.6889, 154.5599, 158.5833, 162.7348, 166.9836, 171.294, 
    175.6264, 179.9403, -175.8037, -171.6418, -167.6047, -163.717, -159.9964, 
    -156.4543, -153.0961, -149.9222, -146.9293, -144.111, -141.459, 
    -138.9637, -136.6147, -134.4015, -132.3136, -130.3409, -128.4736, 
    -126.7026, -125.0193, -123.4158, -121.8846, -120.4189, -119.0124, 
    -117.6592, -116.354, -115.0919, -113.8684, -112.6793, -111.5208, 
    -110.3895, -109.2824, -108.1964, -107.1293, -106.0786, -105.0422, 
    -104.0181, -103.0042, -101.9982, -100.9977, -100, -99.0023, -98.00179, 
    -96.99581, -95.98189, -94.95779, -93.92142, -92.87072, -91.80355, 
    -90.71764, -89.61045, -88.47917, -87.3207, -86.13159, -84.90807, 
    -83.64597, -82.3408, -80.98763, -79.58109, -78.11539, -76.5842, 
    -74.98067, -73.29742, -71.52644, -69.65916, -67.68642, -65.59851, 
    -63.38529, -61.03629, -58.54095, -55.88895, -53.07068, -50.07777, 
    -46.90391, -43.54567, -40.00356, -36.283, -32.39528, -28.3582, -24.19628, 
    -19.94035, -15.62643, -11.29399, -6.983641, -2.734778, 1.416702, 
    5.440118, 9.311138, 13.01213, 16.53197, 19.86536, 23.01188, 25.97502, 
    28.76111, 31.37849, 33.83677, 36.14619, 38.31726, 40.36036, 42.28555, 
    44.10244, 45.82011, 47.44704, 48.99113, 50.45973, 51.85961, 53.19707, 
    54.47794, 55.70762, 56.89116, 58.0333, 59.13849, 60.21099, 61.25488, 
    62.27413, 63.27269, 64.25452, 65.2237, 66.18452, 67.14164, 68.10023, 
    69.06623, 70.04669, 71.05024, 72.08775, 73.17329, 74.32531, 75.56729, 
    76.92528, 78.41363, 80,
  78.44234, 80, 81.55766, 82.98825, 84.26567, 85.41858, 86.48081, 87.47878, 
    88.43163, 89.35334, 90.25443, 91.14309, 92.02596, 92.90859, 93.79587, 
    94.69215, 95.60149, 96.52779, 97.47485, 98.44648, 99.44655, 100.4791, 
    101.5483, 102.6587, 103.8151, 105.0227, 106.2869, 107.614, 109.0107, 
    110.4841, 112.0424, 113.6941, 115.4489, 117.3172, 119.3101, 121.4398, 
    123.719, 126.161, 128.7795, 131.5876, 134.5979, 137.821, 141.2645, 
    144.9315, 148.8196, 152.9183, 157.2088, 161.6623, 166.2411, 170.8996, 
    175.5867, -179.7507, -175.1636, -170.6981, -166.3922, -162.2747, 
    -158.3651, -154.6738, -151.2037, -147.9518, -144.9105, -142.0692, 
    -139.4154, -136.9359, -134.6169, -132.4451, -130.4076, -128.4922, 
    -126.6876, -124.9834, -123.3698, -121.838, -120.38, -118.9885, -117.6567, 
    -116.3785, -115.1485, -113.9616, -112.8132, -111.6993, -110.6162, 
    -109.5605, -108.5295, -107.5205, -106.5315, -105.5604, -104.6054, 
    -103.6649, -102.7368, -101.8186, -100.9075, -100, -99.09254, -98.18142, 
    -97.26324, -96.33508, -95.39455, -94.43964, -93.46854, -92.47948, 
    -91.47052, -90.43948, -89.38383, -88.30069, -87.18678, -86.03842, 
    -84.8515, -83.62148, -82.34333, -81.01153, -79.61997, -78.16199, 
    -76.63023, -75.01662, -73.31236, -71.50779, -69.59242, -67.55492, 
    -65.38312, -63.06414, -60.58459, -57.93084, -55.08951, -52.04818, 
    -48.79626, -45.32621, -41.63491, -37.72529, -33.60784, -29.30191, 
    -24.83636, -20.2493, -15.58666, -10.89963, -6.241157, -1.662304, 
    2.791241, 7.081659, 11.1804, 15.06844, 18.73555, 22.17901, 25.40207, 
    28.41238, 31.22053, 33.83897, 36.281, 38.5602, 40.68988, 42.68283, 
    44.55109, 46.3059, 47.95765, 49.51588, 50.98932, 52.38596, 53.71308, 
    54.97735, 56.18488, 57.34126, 58.45168, 59.52091, 60.55346, 61.55352, 
    62.52515, 63.4722, 64.39851, 65.30785, 66.20413, 67.09141, 67.97404, 
    68.85691, 69.74557, 70.64666, 71.56837, 72.52122, 73.51919, 74.58142, 
    75.73433, 77.01175, 78.44234, 80,
  78.4762, 80, 81.5238, 82.88399, 84.06937, 85.12598, 86.09435, 87.00244, 
    87.8693, 88.70832, 89.52936, 90.34001, 91.14642, 91.95369, 92.76633, 
    93.58841, 94.4237, 95.27586, 96.1485, 97.04527, 97.9699, 98.92633, 
    99.91869, 100.9514, 102.0294, 103.1577, 104.3421, 105.589, 106.9053, 
    108.2986, 109.7776, 111.3516, 113.0314, 114.8284, 116.7557, 118.8273, 
    121.0587, 123.4664, 126.0679, 128.8811, 131.9237, 135.2123, 138.7605, 
    142.5775, 146.6654, 151.0166, 155.612, 160.4184, 165.3891, 170.465, 
    175.5786, -179.3406, -174.3605, -169.5404, -164.9276, -160.5556, 
    -156.4444, -152.6015, -149.0253, -145.7069, -142.6325, -139.7858, 
    -137.1489, -134.7039, -132.4331, -130.32, -128.349, -126.5058, -124.7774, 
    -123.1521, -121.6192, -120.169, -118.793, -117.4834, -116.2332, 
    -115.0362, -113.8867, -112.7797, -111.7106, -110.6755, -109.6709, 
    -108.6936, -107.7413, -106.8117, -105.9032, -105.0144, -104.144, 
    -103.2907, -102.4527, -101.6274, -100.8113, -100, -99.18874, -98.37263, 
    -97.54729, -96.70926, -95.85596, -94.98559, -94.09677, -93.18827, 
    -92.2587, -91.30636, -90.32914, -89.32449, -88.28938, -87.22031, 
    -86.11328, -84.96378, -83.76675, -82.51658, -81.20699, -79.83099, 
    -78.38084, -76.8479, -75.22258, -73.49422, -71.65105, -69.68002, 
    -67.56689, -65.29614, -62.85109, -60.21421, -57.36747, -54.2931, 
    -50.97465, -47.39847, -43.55564, -39.44435, -35.0724, -30.45962, 
    -25.6395, -20.65936, -15.57862, -10.46499, -5.389078, -0.4184048, 
    4.388018, 8.983349, 13.33464, 17.42249, 21.23948, 24.78772, 28.07628, 
    31.11891, 33.9321, 36.53357, 38.94128, 41.17268, 43.24431, 45.17158, 
    46.96864, 48.64837, 50.22244, 51.7014, 53.09473, 54.41098, 55.65785, 
    56.84231, 57.97064, 59.04856, 60.08131, 61.07367, 62.03009, 62.95473, 
    63.8515, 64.72414, 65.5763, 66.41159, 67.23367, 68.04631, 68.85358, 
    69.65999, 70.47064, 71.29168, 72.1307, 72.99756, 73.90565, 74.87402, 
    75.93063, 77.11601, 78.4762, 80,
  78.51732, 80, 81.48268, 82.75737, 83.83998, 84.79482, 85.66682, 86.48399, 
    87.26445, 88.0206, 88.76144, 89.49387, 90.22343, 90.95477, 91.69198, 
    92.43877, 93.19865, 93.97501, 94.77122, 95.59074, 96.43712, 97.31413, 
    98.22578, 99.17644, 100.1708, 101.2141, 102.312, 103.471, 104.6982, 
    106.0015, 107.3899, 108.8736, 110.4639, 112.1737, 114.0174, 116.0114, 
    118.1736, 120.5241, 123.0849, 125.8794, 128.9319, 132.2669, 135.9065, 
    139.8691, 144.165, 148.793, 153.7357, 158.9563, 164.3969, 169.98, 
    175.6142, -178.7972, -173.3458, -168.1098, -163.1479, -158.4976, 
    -154.1769, -150.1875, -146.5193, -143.1543, -140.0701, -137.2426, 
    -134.6471, -132.2601, -130.0597, -128.0256, -126.1396, -124.3852, 
    -122.7479, -121.2148, -119.7741, -118.4159, -117.1309, -115.9112, 
    -114.7496, -113.6397, -112.5759, -111.5532, -110.5672, -109.6141, 
    -108.6906, -107.7941, -106.9224, -106.0739, -105.2477, -104.4432, 
    -103.6597, -102.8967, -102.1527, -101.425, -100.7093, -100, -99.29072, 
    -98.57501, -97.84727, -97.10326, -96.34027, -95.55685, -94.75227, 
    -93.92606, -93.07761, -92.20591, -91.30938, -90.38591, -89.43281, 
    -88.44681, -87.4241, -86.3603, -85.2504, -84.08878, -82.86906, -81.5841, 
    -80.22585, -78.78524, -77.25206, -75.61478, -73.86042, -71.97438, 
    -69.94028, -67.73985, -65.35292, -62.75745, -59.92988, -56.84574, 
    -53.48073, -49.81249, -45.82307, -41.50236, -36.8521, -31.89019, 
    -26.6542, -21.20284, -15.6142, -9.980037, -4.396942, 1.043667, 6.264325, 
    11.20704, 15.83499, 20.13088, 24.09346, 27.73314, 31.06805, 34.1206, 
    36.91507, 39.47586, 41.82642, 43.98864, 45.98256, 47.82631, 49.53611, 
    51.12643, 52.61011, 53.99854, 55.30185, 56.529, 57.68798, 58.78592, 
    59.8292, 60.82357, 61.77421, 62.68587, 63.56288, 64.40926, 65.22878, 
    66.02499, 66.80135, 67.56123, 68.30802, 69.04523, 69.77657, 70.50613, 
    71.23856, 71.9794, 72.73555, 73.51601, 74.33318, 75.20518, 76.16002, 
    77.24263, 78.51732, 80,
  78.56875, 80, 81.43125, 82.60367, 83.5747, 84.4245, 85.19926, 85.92559, 
    86.62003, 87.29374, 87.95471, 88.60906, 89.26173, 89.91685, 90.57809, 
    91.24882, 91.9322, 92.63134, 93.34937, 94.08949, 94.85504, 95.64959, 
    96.47696, 97.34132, 98.24725, 99.19981, 100.2047, 101.2682, 102.3975, 
    103.6006, 104.8869, 106.2668, 107.7524, 109.3574, 111.0977, 112.9914, 
    115.0593, 117.3248, 119.8147, 122.5587, 125.5892, 128.9402, 132.6463, 
    136.7388, 141.2419, 146.1663, 151.502, 157.2107, 163.2212, 169.4302, 
    175.7105, -178.0743, -172.052, -166.3267, -160.9707, -156.0232, 
    -151.4949, -147.3757, -143.6418, -140.2616, -137.2009, -134.4254, 
    -131.9025, -129.6025, -127.4984, -125.5666, -123.7862, -122.1388, 
    -120.6084, -119.1812, -117.845, -116.5891, -115.4043, -114.2822, 
    -113.2159, -112.1989, -111.2256, -110.2914, -109.3918, -108.5234, 
    -107.6833, -106.8691, -106.0792, -105.3128, -104.5698, -103.8505, 
    -103.1556, -102.4853, -101.8385, -101.2125, -100.6021, -100, -99.39791, 
    -98.78746, -98.16146, -97.51475, -96.84442, -96.14951, -95.43023, 
    -94.68719, -93.92081, -93.13094, -92.31672, -91.47656, -90.60818, 
    -89.70864, -88.77436, -87.80114, -86.78412, -85.71776, -84.59574, 
    -83.41087, -82.15499, -80.81876, -79.39157, -77.86124, -76.21383, 
    -74.43337, -72.50157, -70.39754, -68.0975, -65.57463, -62.7991, -59.7384, 
    -56.35823, -52.62425, -48.50509, -43.97684, -39.02929, -33.67328, 
    -27.94805, -21.92572, -15.71052, -9.43022, -3.221188, 2.789308, 8.497978, 
    13.83367, 18.75813, 23.26125, 27.35374, 31.05976, 34.41084, 37.44126, 
    40.18525, 42.67518, 44.94074, 47.00857, 48.90226, 50.64256, 52.24758, 
    53.73316, 55.11308, 56.39937, 57.60255, 58.73183, 59.79533, 60.80019, 
    61.75275, 62.65868, 63.52304, 64.35041, 65.14496, 65.91051, 66.65063, 
    67.36866, 68.0678, 68.75118, 69.42191, 70.08315, 70.73827, 71.39094, 
    72.04529, 72.70626, 73.37997, 74.07441, 74.80074, 75.5755, 76.4253, 
    77.39633, 78.56875, 80,
  78.63466, 80, 81.36534, 82.41873, 83.27239, 84.01614, 84.69427, 85.33079, 
    85.94028, 86.53245, 87.11426, 87.69102, 88.26704, 88.84595, 89.43098, 
    90.02511, 90.63118, 91.252, 91.8904, 92.5493, 93.2318, 93.9412, 94.68106, 
    95.45531, 96.2683, 97.12486, 98.03043, 98.99117, 100.0141, 101.1072, 
    102.2797, 103.5423, 104.9073, 106.3891, 108.0044, 109.7729, 111.7177, 
    113.8654, 116.2476, 118.9003, 121.865, 125.1877, 128.9184, 133.1074, 
    137.8006, 143.0303, 148.8036, 155.0875, 161.7974, 168.7936, 175.8931, 
    -177.1043, -170.3822, -164.0817, -158.2885, -153.0367, -148.32, 
    -144.1064, -140.3502, -137.0009, -134.0088, -131.3274, -128.9152, 
    -126.7358, -124.7577, -122.9539, -121.3012, -119.7798, -118.3728, 
    -117.0656, -115.8458, -114.7026, -113.6266, -112.6098, -111.6451, 
    -110.7263, -109.8481, -109.0059, -108.1957, -107.4143, -106.659, 
    -105.928, -105.2204, -104.5361, -103.8761, -103.2422, -102.6364, 
    -102.0602, -101.5133, -100.9923, -100.4909, -100, -99.50912, -99.00771, 
    -98.48674, -97.93977, -97.36359, -96.75783, -96.12391, -95.46393, 
    -94.77965, -94.07203, -93.34105, -92.58574, -91.80428, -90.99409, 
    -90.15188, -89.2737, -88.35492, -87.3902, -86.37337, -85.2974, -84.15417, 
    -82.93436, -81.6272, -80.22018, -78.6988, -77.0461, -75.24228, -73.26421, 
    -71.08482, -68.67262, -65.99121, -62.99907, -59.64984, -55.89364, -51.68, 
    -46.96329, -41.71145, -35.91832, -29.61777, -22.89572, -15.89308, 
    -8.793619, -1.797381, 4.912534, 11.19644, 16.96969, 22.19945, 26.8926, 
    31.08161, 34.81226, 38.13502, 41.09968, 43.75241, 46.13455, 48.28233, 
    50.22705, 51.9956, 53.61095, 55.09272, 56.45771, 57.72029, 58.89281, 
    59.98592, 61.00883, 61.96957, 62.87514, 63.7317, 64.54469, 65.31894, 
    66.0588, 66.7682, 67.4507, 68.1096, 68.748, 69.36882, 69.97489, 70.56902, 
    71.15405, 71.73296, 72.30898, 72.88574, 73.46755, 74.05972, 74.66921, 
    75.30573, 75.98386, 76.72761, 77.58127, 78.63466, 80,
  78.72022, 80, 81.27978, 82.1999, 82.93392, 83.57271, 84.15597, 84.70443, 
    85.23051, 85.74244, 86.24611, 86.74606, 87.24596, 87.74892, 88.25777, 
    88.77508, 89.30335, 89.84507, 90.40275, 90.97902, 91.57666, 92.19866, 
    92.8483, 93.52915, 94.24524, 95.00107, 95.80174, 96.65305, 97.56169, 
    98.53534, 99.58294, 100.7149, 101.9436, 103.2834, 104.7516, 106.3685, 
    108.1588, 110.1518, 112.3829, 114.8944, 117.7367, 120.9693, 124.6607, 
    128.8866, 133.7249, 139.2451, 145.4897, 152.4476, 160.0265, 168.0358, 
    176.2016, -175.7835, -168.1943, -161.2224, -154.9615, -149.4234, 
    -144.5661, -140.3203, -136.6081, -133.3535, -130.4881, -127.9522, 
    -125.695, -123.6742, -121.8542, -120.2055, -118.7034, -117.3273, 
    -116.0598, -114.8864, -113.7945, -112.7737, -111.8149, -110.9102, 
    -110.0529, -109.2372, -108.458, -107.7111, -106.9926, -106.2998, 
    -105.6302, -104.9827, -104.3569, -103.7538, -103.1757, -102.6262, 
    -102.1092, -101.6279, -101.1822, -100.7683, -100.3779, -100, -99.62212, 
    -99.23173, -98.81776, -98.37212, -97.89077, -97.37383, -96.8243, 
    -96.24619, -95.64307, -95.01727, -94.36977, -93.70025, -93.00739, 
    -92.28895, -91.54197, -90.76279, -89.9471, -89.08983, -88.18513, 
    -87.2263, -86.20548, -85.11364, -83.94019, -82.67271, -81.29659, 
    -79.79449, -78.14578, -76.32579, -74.30497, -72.04783, -69.51187, 
    -66.64645, -63.39194, -59.67973, -55.43391, -50.57658, -45.03846, 
    -38.77757, -31.80567, -24.21651, -16.20164, -8.035747, -0.02645781, 
    7.55235, 14.51032, 20.75487, 26.2751, 31.11345, 35.33934, 39.0307, 
    42.26331, 45.10563, 47.61708, 49.84815, 51.84118, 53.63147, 55.24844, 
    56.71658, 58.05639, 59.28506, 60.41706, 61.46466, 62.43831, 63.34694, 
    64.19826, 64.99893, 65.75476, 66.47085, 67.1517, 67.80134, 68.42334, 
    69.02098, 69.59725, 70.15493, 70.69665, 71.22492, 71.74223, 72.25108, 
    72.75404, 73.25394, 73.75389, 74.25756, 74.76949, 75.29557, 75.84403, 
    76.42729, 77.06608, 77.8001, 78.72022, 80,
  78.83092, 80, 81.16908, 81.94684, 82.56233, 83.0988, 83.58978, 84.05244, 
    84.49699, 84.93024, 85.35705, 85.78119, 86.20573, 86.63329, 87.06626, 
    87.50684, 87.95717, 88.41939, 88.89568, 89.38835, 89.89982, 90.43274, 
    90.99001, 91.57481, 92.19077, 92.84193, 93.53293, 94.26905, 95.05643, 
    95.90222, 96.81477, 97.80392, 98.88142, 100.0612, 101.3603, 102.799, 
    104.4023, 106.201, 108.2328, 110.5448, 113.1954, 116.2568, 119.8177, 
    123.9844, 128.8792, 134.63, 141.3473, 149.079, 157.7484, 167.099, 
    176.702, -173.9455, -165.2725, -157.5354, -150.8111, -145.0516, 
    -140.1466, -135.9678, -132.3932, -129.3163, -126.6485, -124.3172, 
    -122.2642, -120.4422, -118.8134, -117.347, -116.0179, -114.8055, 
    -113.6929, -112.6658, -111.7125, -110.823, -109.9886, -109.2022, 
    -108.4575, -107.7491, -107.0724, -106.4234, -105.7986, -105.1956, 
    -104.6123, -104.0479, -103.5027, -102.9787, -102.4802, -102.0131, 
    -101.584, -101.1977, -100.8542, -100.5474, -100.267, -100, -99.73305, 
    -99.45258, -99.14581, -98.80226, -98.41599, -97.98692, -97.51979, 
    -97.02126, -96.49734, -95.95215, -95.38772, -94.80444, -94.20138, 
    -93.57664, -92.92759, -92.25085, -91.54247, -90.79778, -90.01139, 
    -89.17705, -88.28748, -87.33417, -86.30711, -85.19447, -83.98209, 
    -82.65298, -81.18657, -79.55779, -77.73585, -75.68279, -73.35153, 
    -70.68365, -67.60679, -64.03219, -59.85344, -54.9484, -49.18893, 
    -42.46464, -34.7275, -26.05452, -16.702, -7.099045, 2.251643, 10.92097, 
    18.65274, 25.37001, 31.12083, 36.01556, 40.18235, 43.74324, 46.80462, 
    49.45517, 51.76719, 53.79903, 55.59768, 57.20101, 58.63971, 59.93876, 
    61.11859, 62.19608, 63.18523, 64.09778, 64.94357, 65.73095, 66.46707, 
    67.15807, 67.80923, 68.42519, 69.00999, 69.56726, 70.10018, 70.61165, 
    71.10432, 71.58061, 72.04283, 72.49316, 72.93374, 73.36671, 73.79427, 
    74.21881, 74.64295, 75.06976, 75.50301, 75.94756, 76.41022, 76.9012, 
    77.43767, 78.05316, 78.83092, 80,
  78.97098, 80, 81.02902, 81.66203, 82.16265, 82.60043, 83.00219, 83.38155, 
    83.74667, 84.10297, 84.45437, 84.80391, 85.15408, 85.50705, 85.86475, 
    86.229, 86.6016, 86.98433, 87.37902, 87.78761, 88.21217, 88.65494, 
    89.11839, 89.60529, 90.11873, 90.66222, 91.23981, 91.85614, 92.51659, 
    93.22752, 93.99638, 94.83207, 95.74525, 96.74881, 97.85847, 99.09361, 
    100.4783, 102.0426, 103.825, 105.8741, 108.2533, 111.0442, 114.3537, 
    118.3198, 123.118, 128.9603, 136.0754, 144.6475, 154.6891, 165.8801, 
    177.5113, -171.3072, -161.2801, -152.7229, -145.6194, -139.7845, 
    -134.9892, -131.022, -127.7078, -124.909, -122.5191, -120.4564, 
    -118.6581, -117.0753, -115.6697, -114.4112, -113.2756, -112.2436, 
    -111.2994, -110.4298, -109.6242, -108.8734, -108.1698, -107.5069, 
    -106.8792, -106.2817, -105.7103, -105.1615, -104.6321, -104.1198, 
    -103.6229, -103.1407, -102.6741, -102.2264, -101.804, -101.4167, 
    -101.0749, -100.7847, -100.5435, -100.3411, -100.1644, -100, -99.83563, 
    -99.65885, -99.4565, -99.21532, -98.92513, -98.58331, -98.19596, 
    -97.77359, -97.32589, -96.85931, -96.37711, -95.88017, -95.36787, 
    -94.83852, -94.28968, -93.71832, -93.12085, -92.4931, -91.83022, 
    -91.12665, -90.37585, -89.57019, -88.70063, -87.75636, -86.72437, 
    -85.58883, -84.33032, -82.92474, -81.34189, -79.54356, -77.48092, 
    -75.09102, -72.29217, -68.97798, -65.01076, -60.21552, -54.38064, 
    -47.27715, -38.71988, -28.69284, -17.51129, -5.880136, 5.310857, 
    15.35251, 23.92456, 31.03975, 36.88199, 41.68015, 45.64628, 48.95577, 
    51.74675, 54.12586, 56.17503, 57.95735, 59.52172, 60.90639, 62.14153, 
    63.25119, 64.25475, 65.16793, 66.00362, 66.77248, 67.48341, 68.14386, 
    68.76019, 69.33778, 69.88127, 70.39471, 70.88161, 71.34506, 71.78783, 
    72.21239, 72.62098, 73.01567, 73.3984, 73.771, 74.13525, 74.49295, 
    74.84592, 75.19609, 75.54563, 75.89703, 76.25333, 76.61845, 76.99781, 
    77.39957, 77.83735, 78.33797, 78.97098, 80,
  79.14133, 80, 80.85867, 81.35062, 81.7415, 82.08465, 82.40038, 82.69906, 
    82.98692, 83.26811, 83.5457, 83.82202, 84.09904, 84.37843, 84.66174, 
    84.95042, 85.24588, 85.54954, 85.86289, 86.18747, 86.52497, 86.87719, 
    87.24616, 87.63412, 88.04362, 88.47755, 88.93924, 89.43253, 89.96194, 
    90.53278, 91.15134, 91.82516, 92.56339, 93.37716, 94.28021, 95.28966, 
    96.42711, 97.72015, 99.20451, 100.9271, 102.9506, 105.3598, 108.2711, 
    111.8468, 116.3132, 121.9823, 129.2628, 138.6142, 150.3448, 164.1736, 
    178.8606, -167.3524, -155.6814, -146.3857, -139.148, -133.5086, 
    -129.0614, -125.4965, -122.5896, -120.1799, -118.1518, -116.4212, 
    -114.9258, -113.6189, -112.465, -111.4366, -110.5121, -109.6743, 
    -108.9095, -108.2063, -107.5556, -106.9496, -106.3817, -105.8466, 
    -105.3393, -104.8558, -104.3924, -103.9459, -103.5136, -103.0931, 
    -102.6827, -102.2817, -101.8912, -101.5155, -101.1647, -100.8554, 
    -100.604, -100.4142, -100.2743, -100.1675, -100.0795, -100, -99.92047, 
    -99.83251, -99.72566, -99.58578, -99.39602, -99.14462, -98.83527, 
    -98.48452, -98.10884, -97.71828, -97.31728, -96.9069, -96.4864, 
    -96.05408, -95.6076, -95.1442, -94.66068, -94.15342, -93.61826, 
    -93.05044, -92.44441, -91.79369, -91.09054, -90.32569, -89.48792, 
    -88.5634, -87.535, -86.38111, -85.07424, -83.57882, -81.84816, -79.82008, 
    -77.41041, -74.5035, -70.93864, -66.49138, -60.85201, -53.61435, 
    -44.31855, -32.64756, -18.86065, -4.173635, 9.655166, 21.38583, 30.7372, 
    38.01767, 43.68684, 48.15319, 51.72887, 54.64023, 57.04939, 59.07287, 
    60.79549, 62.27985, 63.57289, 64.71034, 65.71979, 66.62284, 67.43661, 
    68.17484, 68.84866, 69.46722, 70.03806, 70.56747, 71.06076, 71.52245, 
    71.95638, 72.36588, 72.75384, 73.12281, 73.47503, 73.81253, 74.13711, 
    74.45046, 74.75412, 75.04958, 75.33826, 75.62157, 75.90096, 76.17798, 
    76.4543, 76.73189, 77.01308, 77.30094, 77.59962, 77.91535, 78.2585, 
    78.64938, 79.14133, 80,
  79.33845, 80, 80.66155, 81.01993, 81.30656, 81.55907, 81.79189, 82.01244, 
    82.2252, 82.43322, 82.63869, 82.84333, 83.04858, 83.25569, 83.46578, 
    83.67994, 83.89921, 84.12466, 84.35741, 84.5986, 84.84952, 85.11151, 
    85.38612, 85.67503, 85.9802, 86.30383, 86.64845, 87.01702, 87.41303, 
    87.84057, 88.30454, 88.81084, 89.36665, 89.98077, 90.66421, 91.43075, 
    92.29802, 93.28888, 94.43342, 95.77206, 97.36021, 99.27563, 101.6303, 
    104.5898, 108.4062, 113.4719, 120.402, 130.1146, 143.707, 161.5079, 
    -178.7233, -161.0628, -147.6345, -138.0468, -131.1994, -126.1864, 
    -122.4029, -119.4634, -117.1198, -115.2091, -113.6209, -112.2785, 
    -111.127, -110.1264, -109.2469, -108.4658, -107.7654, -107.1321, 
    -106.5547, -106.0243, -105.5337, -105.0768, -104.6484, -104.2441, 
    -103.8602, -103.4932, -103.1403, -102.7985, -102.4654, -102.1385, 
    -101.8157, -101.4954, -101.1777, -100.8678, -100.5836, -100.3603, 
    -100.2179, -100.1355, -100.0851, -100.0506, -100.0237, -100, -99.97626, 
    -99.94939, -99.91489, -99.86455, -99.78211, -99.63968, -99.41637, 
    -99.13221, -98.82231, -98.50465, -98.18433, -97.8615, -97.5346, 
    -97.20148, -96.85972, -96.50676, -96.13983, -95.75591, -95.35165, 
    -94.92323, -94.46629, -93.97568, -93.44534, -92.86794, -92.2346, 
    -91.53424, -90.75311, -89.8736, -88.87302, -87.7215, -86.37905, 
    -84.79086, -82.88018, -80.53661, -77.59708, -73.81362, -68.80055, 
    -61.95322, -52.36549, -38.93719, -21.2767, -1.507927, 16.29298, 29.88544, 
    39.59801, 46.52807, 51.59385, 55.41024, 58.36973, 60.72436, 62.63979, 
    64.22794, 65.56658, 66.71112, 67.70198, 68.56925, 69.33579, 70.01923, 
    70.63335, 71.18916, 71.69546, 72.15943, 72.58697, 72.98298, 73.35155, 
    73.69617, 74.0198, 74.32497, 74.61388, 74.88849, 75.15048, 75.4014, 
    75.64259, 75.87534, 76.10079, 76.32006, 76.53422, 76.74431, 76.95142, 
    77.15667, 77.36131, 77.56678, 77.7748, 77.98756, 78.20811, 78.44093, 
    78.69344, 78.98007, 79.33845, 80,
  79.55453, 80, 80.44547, 80.67855, 80.86597, 81.03147, 81.18425, 81.3291, 
    81.46893, 81.60568, 81.74081, 81.87543, 82.01049, 82.1468, 82.28511, 
    82.42612, 82.57053, 82.71906, 82.87241, 83.03138, 83.19679, 83.36958, 
    83.55073, 83.7414, 83.94289, 84.15666, 84.38444, 84.6282, 84.8903, 
    85.17352, 85.48118, 85.8173, 86.1868, 86.59574, 87.05174, 87.5644, 
    88.14613, 88.81317, 89.58716, 90.49764, 91.58596, 92.91167, 94.56358, 
    96.67969, 99.48489, 103.3674, 109.041, 117.8948, 132.5935, 156.5226, 
    -173.7402, -150.2899, -135.9617, -127.3108, -121.7468, -117.9264, 
    -115.1577, -113.0634, -111.424, -110.1047, -109.0184, -108.1066, 
    -107.3286, -106.6552, -106.0651, -105.5422, -105.0742, -104.6513, 
    -104.2661, -103.9122, -103.5848, -103.2795, -102.9929, -102.7218, 
    -102.4636, -102.2158, -101.9761, -101.7423, -101.5119, -101.2823, 
    -101.0504, -100.8122, -100.563, -100.3058, -100.1113, -100.0426, 
    -100.0209, -100.0119, -100.007, -100.0041, -100.0019, -100, -99.99806, 
    -99.99586, -99.99296, -99.98814, -99.97906, -99.9574, -99.88869, 
    -99.69417, -99.43704, -99.18782, -98.94959, -98.7177, -98.48813, 
    -98.25772, -98.02386, -97.78416, -97.53637, -97.27818, -97.00711, 
    -96.72048, -96.41522, -96.08775, -95.73392, -95.34866, -94.92581, 
    -94.45776, -93.93486, -93.34479, -92.67145, -91.89345, -90.98164, 
    -89.8953, -88.57598, -86.93661, -84.84226, -82.07361, -78.2532, 
    -72.68923, -64.03826, -49.71014, -26.25977, 3.477372, 27.40649, 42.10522, 
    50.95898, 56.63261, 60.51511, 63.32031, 65.43642, 67.08833, 68.41404, 
    69.50236, 70.41284, 71.18683, 71.85387, 72.4356, 72.94826, 73.40426, 
    73.8132, 74.1827, 74.51882, 74.82648, 75.1097, 75.3718, 75.61556, 
    75.84334, 76.05711, 76.2586, 76.44927, 76.63042, 76.80321, 76.96862, 
    77.12759, 77.28094, 77.42947, 77.57388, 77.71489, 77.8532, 77.98951, 
    78.12457, 78.25919, 78.39432, 78.53107, 78.6709, 78.81575, 78.96853, 
    79.13403, 79.32145, 79.55453, 80,
  79.77896, 80, 80.22104, 80.33562, 80.4279, 80.50944, 80.58473, 80.65613, 
    80.72506, 80.79248, 80.8591, 80.92548, 80.99207, 81.05929, 81.12749, 
    81.19703, 81.26825, 81.3415, 81.41714, 81.49555, 81.57716, 81.6624, 
    81.75179, 81.84589, 81.94534, 82.0509, 82.16338, 82.28381, 82.41333, 
    82.55336, 82.70555, 82.87193, 83.05496, 83.25774, 83.48408, 83.73889, 
    84.02854, 84.36134, 84.74855, 85.20562, 85.75446, 86.42712, 87.2725, 
    88.36884, 89.84963, 91.96172, 95.21452, 100.8343, 112.489, 143.331, 
    -159.9273, -130.8179, -119.7029, -114.2738, -111.1055, -109.0369, 
    -107.5803, -106.498, -105.6607, -104.9923, -104.4451, -103.9876, 
    -103.5984, -103.2623, -102.9682, -102.7079, -102.4749, -102.2645, 
    -102.0727, -101.8964, -101.7331, -101.5806, -101.437, -101.3008, 
    -101.1706, -101.0448, -100.9221, -100.8011, -100.6798, -100.5557, 
    -100.4245, -100.2761, -100.071, -100.0002, -100.0001, -100.0001, 
    -100.0001, -100.0001, -100.0001, -100, -100, -100, -99.99998, -99.99996, 
    -99.99995, -99.99992, -99.99991, -99.99989, -99.99987, -99.99985, 
    -99.92899, -99.72395, -99.57553, -99.44427, -99.32018, -99.19891, 
    -99.07788, -98.95522, -98.82944, -98.69916, -98.56297, -98.4194, 
    -98.26688, -98.10355, -97.92728, -97.7355, -97.52507, -97.29213, 
    -97.03176, -96.73766, -96.40156, -96.01239, -95.55492, -95.00766, 
    -94.33926, -93.50198, -92.4197, -90.96311, -88.89446, -85.72624, 
    -80.29715, -69.18208, -40.07274, 16.66903, 47.51101, 59.16573, 64.78548, 
    68.03828, 70.15037, 71.63116, 72.7275, 73.57288, 74.24554, 74.79438, 
    75.25145, 75.63866, 75.97146, 76.26111, 76.51592, 76.74226, 76.94504, 
    77.12807, 77.29445, 77.44664, 77.58667, 77.71619, 77.83662, 77.9491, 
    78.05466, 78.15411, 78.24821, 78.3376, 78.42284, 78.50445, 78.58286, 
    78.6585, 78.73175, 78.80297, 78.87251, 78.94071, 79.00793, 79.07452, 
    79.1409, 79.20752, 79.27494, 79.34387, 79.41527, 79.49056, 79.5721, 
    79.66438, 79.77896, 80,
  80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 
    80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 
    80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, -100, -100, -100, 
    -100, -100, -100, -100, -100, -100, -100, -100, -100, -100, -100, -100, 
    -100, -100, -100, -100, -100, -100, -100, -100, -100, -100, -100, -100, 
    -100, -100, -100, -100, -100, -100, -100, -100, -100, -100, -100, -100, 
    -100, -100, -100, -100, -100, -100, -100, -100, -100, -100, -100, -100, 
    -100, -100, -100, -100, -100, -100, -100, -100, -100, -100, -100, -100, 
    -100, -100, -100, -100, -100, -100, -100, -100, -100, -100, -100, -100, 
    -100, -100, -100, -100, -100, -100, -100, -100, 80, 80, 80, 80, 80, 80, 
    80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 
    80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 
    80, 80, 80, 80, 80, 80, 80,
  80.22104, 80, 79.77896, 79.66438, 79.5721, 79.49056, 79.41527, 79.34387, 
    79.27494, 79.20752, 79.1409, 79.07452, 79.00793, 78.94071, 78.87251, 
    78.80297, 78.73175, 78.6585, 78.58286, 78.50445, 78.42284, 78.3376, 
    78.24821, 78.15411, 78.05466, 77.9491, 77.83662, 77.71619, 77.58667, 
    77.44664, 77.29445, 77.12807, 76.94504, 76.74226, 76.51592, 76.26111, 
    75.97146, 75.63866, 75.25145, 74.79438, 74.24554, 73.57288, 72.7275, 
    71.63116, 70.15037, 68.03828, 64.78548, 59.16573, 47.51101, 16.66903, 
    -40.07274, -69.18208, -80.29715, -85.72624, -88.89446, -90.96311, 
    -92.4197, -93.50198, -94.33926, -95.00766, -95.55492, -96.01239, 
    -96.40156, -96.73766, -97.03176, -97.29213, -97.52507, -97.7355, 
    -97.92728, -98.10355, -98.26688, -98.4194, -98.56297, -98.69916, 
    -98.82944, -98.95522, -99.07788, -99.19891, -99.32018, -99.44427, 
    -99.57553, -99.72395, -99.92899, -99.99985, -99.99987, -99.99989, 
    -99.99991, -99.99992, -99.99995, -99.99996, -99.99998, -100, -100, -100, 
    -100.0001, -100.0001, -100.0001, -100.0001, -100.0001, -100.0002, 
    -100.071, -100.2761, -100.4245, -100.5557, -100.6798, -100.8011, 
    -100.9221, -101.0448, -101.1706, -101.3008, -101.437, -101.5806, 
    -101.7331, -101.8964, -102.0727, -102.2645, -102.4749, -102.7079, 
    -102.9682, -103.2623, -103.5984, -103.9876, -104.4451, -104.9923, 
    -105.6607, -106.498, -107.5803, -109.0369, -111.1055, -114.2738, 
    -119.7029, -130.8179, -159.9273, 143.331, 112.489, 100.8343, 95.21452, 
    91.96172, 89.84963, 88.36884, 87.2725, 86.42712, 85.75446, 85.20562, 
    84.74855, 84.36134, 84.02854, 83.73889, 83.48408, 83.25774, 83.05496, 
    82.87193, 82.70555, 82.55336, 82.41333, 82.28381, 82.16338, 82.0509, 
    81.94534, 81.84589, 81.75179, 81.6624, 81.57716, 81.49555, 81.41714, 
    81.3415, 81.26825, 81.19703, 81.12749, 81.05929, 80.99207, 80.92548, 
    80.8591, 80.79248, 80.72506, 80.65613, 80.58473, 80.50944, 80.4279, 
    80.33562, 80.22104, 80 ;

 sic_tot_var =
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5,
  0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5 ;
}
